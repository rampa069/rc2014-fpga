
--
-- Copyright (c) 2008-2023 Sytse van Slooten
--
-- Permission is hereby granted to any person obtaining a copy of these VHDL source files and
-- other language source files and associated documentation files ("the materials") to use
-- these materials solely for personal, non-commercial purposes.
-- You are also granted permission to make changes to the materials, on the condition that this
-- copyright notice is retained unchanged.
--
-- The materials are distributed in the hope that they will be useful, but WITHOUT ANY WARRANTY;
-- without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.
--

-- $Revision$

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity vtbr is
   port(
      base_addr : in std_logic_vector(17 downto 0);

      bus_addr_match : out std_logic;
      bus_addr : in std_logic_vector(17 downto 0);
      bus_dati : out std_logic_vector(15 downto 0);
      bus_dato : in std_logic_vector(15 downto 0);
      bus_control_dati : in std_logic;
      bus_control_dato : in std_logic;
      bus_control_datob : in std_logic;

      reset : in std_logic;
      clk : in std_logic
   );
end vtbr;

architecture implementation of vtbr is

signal base_addr_match : std_logic;

subtype u is std_logic_vector(7 downto 0);
type mem_type is array(0 to 4095) of u;

-- INSERT MEMORY CONTENTS HERE

-- code base at 0

signal meme : mem_type := mem_type'(
u'(x"77"),u'(x"fc"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"01"),u'(x"18"),
u'(x"18"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"01"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"01"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"01"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"01"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"01"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"01"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"01"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"01"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"01"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"df"),u'(x"e0"),u'(x"fe"),u'(x"c6"),u'(x"00"),u'(x"37"),u'(x"d6"),u'(x"37"),u'(x"d4"),u'(x"37"),u'(x"ca"),u'(x"37"),u'(x"c8"),u'(x"37"),u'(x"c5"),u'(x"37"),
u'(x"c6"),u'(x"37"),u'(x"c4"),u'(x"df"),u'(x"b4"),u'(x"30"),u'(x"df"),u'(x"e0"),u'(x"32"),u'(x"df"),u'(x"16"),u'(x"34"),u'(x"df"),u'(x"e0"),u'(x"36"),u'(x"df"),
u'(x"18"),u'(x"38"),u'(x"df"),u'(x"e0"),u'(x"3a"),u'(x"df"),u'(x"40"),u'(x"70"),u'(x"df"),u'(x"40"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"37"),u'(x"24"),
u'(x"f7"),u'(x"26"),u'(x"c3"),u'(x"00"),u'(x"d3"),u'(x"20"),u'(x"d7"),u'(x"00"),u'(x"fb"),u'(x"c2"),u'(x"52"),u'(x"c3"),u'(x"00"),u'(x"df"),u'(x"69"),u'(x"0a"),
u'(x"02"),u'(x"c2"),u'(x"70"),u'(x"80"),u'(x"13"),u'(x"fd"),u'(x"e3"),u'(x"20"),u'(x"37"),u'(x"be"),u'(x"37"),u'(x"bb"),u'(x"37"),u'(x"b8"),u'(x"37"),u'(x"b5"),
u'(x"37"),u'(x"b2"),u'(x"37"),u'(x"af"),u'(x"37"),u'(x"ac"),u'(x"f7"),u'(x"a0"),u'(x"f7"),u'(x"03"),u'(x"36"),u'(x"f7"),u'(x"01"),u'(x"34"),u'(x"f7"),u'(x"01"),
u'(x"2c"),u'(x"f7"),u'(x"01"),u'(x"2a"),u'(x"f7"),u'(x"42"),u'(x"2c"),u'(x"f7"),u'(x"42"),u'(x"24"),u'(x"f7"),u'(x"42"),u'(x"1f"),u'(x"f7"),u'(x"42"),u'(x"1b"),
u'(x"f7"),u'(x"01"),u'(x"16"),u'(x"f7"),u'(x"18"),u'(x"12"),u'(x"f7"),u'(x"18"),u'(x"0e"),u'(x"37"),u'(x"00"),u'(x"37"),u'(x"fd"),u'(x"37"),u'(x"6c"),u'(x"f7"),
u'(x"01"),u'(x"62"),u'(x"37"),u'(x"5d"),u'(x"37"),u'(x"58"),u'(x"37"),u'(x"59"),u'(x"37"),u'(x"53"),u'(x"37"),u'(x"dc"),u'(x"37"),u'(x"d9"),u'(x"37"),u'(x"3b"),
u'(x"37"),u'(x"38"),u'(x"37"),u'(x"31"),u'(x"37"),u'(x"2e"),u'(x"37"),u'(x"38"),u'(x"1f"),u'(x"02"),u'(x"1f"),u'(x"04"),u'(x"1f"),u'(x"06"),u'(x"1f"),u'(x"0c"),
u'(x"f7"),u'(x"e6"),u'(x"1f"),u'(x"00"),u'(x"f7"),u'(x"78"),u'(x"c0"),u'(x"10"),u'(x"9f"),u'(x"0c"),u'(x"f7"),u'(x"32"),u'(x"c0"),u'(x"0a"),u'(x"57"),u'(x"e0"),
u'(x"03"),u'(x"f7"),u'(x"3e"),u'(x"ec"),u'(x"40"),u'(x"f7"),u'(x"9c"),u'(x"e8"),u'(x"f7"),u'(x"f6"),u'(x"c0"),u'(x"e4"),u'(x"9f"),u'(x"0d"),u'(x"c1"),u'(x"80"),
u'(x"f7"),u'(x"94"),u'(x"c1"),u'(x"dc"),u'(x"40"),u'(x"ae"),u'(x"c0"),u'(x"02"),u'(x"37"),u'(x"f0"),u'(x"c0"),u'(x"ec"),u'(x"c0"),u'(x"f1"),u'(x"c0"),u'(x"8e"),
u'(x"00"),u'(x"c8"),u'(x"cd"),u'(x"57"),u'(x"40"),u'(x"0d"),u'(x"57"),u'(x"4c"),u'(x"0a"),u'(x"c1"),u'(x"40"),u'(x"c1"),u'(x"41"),u'(x"26"),u'(x"77"),u'(x"9e"),
u'(x"37"),u'(x"9c"),u'(x"2e"),u'(x"57"),u'(x"20"),u'(x"28"),u'(x"57"),u'(x"3f"),u'(x"25"),u'(x"f7"),u'(x"8a"),u'(x"0d"),u'(x"77"),u'(x"84"),u'(x"c0"),u'(x"7e"),
u'(x"17"),u'(x"58"),u'(x"04"),u'(x"17"),u'(x"b4"),u'(x"01"),u'(x"1a"),u'(x"c8"),u'(x"18"),u'(x"c1"),u'(x"e0"),u'(x"c1"),u'(x"c1"),u'(x"c1"),u'(x"c1"),u'(x"c1"),
u'(x"f7"),u'(x"e0"),u'(x"5a"),u'(x"c1"),u'(x"56"),u'(x"37"),u'(x"52"),u'(x"f7"),u'(x"4c"),u'(x"04"),u'(x"c0"),u'(x"46"),u'(x"c8"),u'(x"03"),u'(x"37"),u'(x"40"),
u'(x"87"),u'(x"00"),u'(x"87"),u'(x"40"),u'(x"58"),u'(x"26"),u'(x"50"),u'(x"7c"),u'(x"a8"),u'(x"a8"),u'(x"a8"),u'(x"aa"),u'(x"b4"),u'(x"2a"),u'(x"4c"),u'(x"78"),
u'(x"c1"),u'(x"00"),u'(x"f7"),u'(x"14"),u'(x"03"),u'(x"5f"),u'(x"04"),u'(x"03"),u'(x"5f"),u'(x"06"),u'(x"00"),u'(x"87"),u'(x"c1"),u'(x"01"),u'(x"04"),u'(x"df"),
u'(x"01"),u'(x"02"),u'(x"03"),u'(x"df"),u'(x"01"),u'(x"02"),u'(x"c1"),u'(x"02"),u'(x"04"),u'(x"df"),u'(x"02"),u'(x"02"),u'(x"03"),u'(x"df"),u'(x"02"),u'(x"02"),
u'(x"c1"),u'(x"04"),u'(x"04"),u'(x"df"),u'(x"04"),u'(x"02"),u'(x"03"),u'(x"df"),u'(x"04"),u'(x"02"),u'(x"c1"),u'(x"08"),u'(x"04"),u'(x"df"),u'(x"08"),u'(x"02"),
u'(x"03"),u'(x"df"),u'(x"08"),u'(x"02"),u'(x"c1"),u'(x"10"),u'(x"04"),u'(x"df"),u'(x"10"),u'(x"02"),u'(x"03"),u'(x"df"),u'(x"10"),u'(x"02"),u'(x"c1"),u'(x"40"),
u'(x"04"),u'(x"df"),u'(x"00"),u'(x"02"),u'(x"03"),u'(x"df"),u'(x"00"),u'(x"02"),u'(x"f7"),u'(x"8c"),u'(x"27"),u'(x"c1"),u'(x"80"),u'(x"04"),u'(x"df"),u'(x"00"),
u'(x"02"),u'(x"03"),u'(x"df"),u'(x"00"),u'(x"02"),u'(x"c1"),u'(x"20"),u'(x"04"),u'(x"f7"),u'(x"01"),u'(x"66"),u'(x"02"),u'(x"37"),u'(x"60"),u'(x"c1"),u'(x"00"),
u'(x"04"),u'(x"df"),u'(x"00"),u'(x"02"),u'(x"03"),u'(x"df"),u'(x"00"),u'(x"02"),u'(x"c1"),u'(x"00"),u'(x"04"),u'(x"df"),u'(x"00"),u'(x"02"),u'(x"03"),u'(x"df"),
u'(x"00"),u'(x"02"),u'(x"87"),u'(x"c0"),u'(x"38"),u'(x"c0"),u'(x"c0"),u'(x"00"),u'(x"c0"),u'(x"00"),u'(x"48"),u'(x"df"),u'(x"00"),u'(x"02"),u'(x"08"),u'(x"b7"),
u'(x"20"),u'(x"f7"),u'(x"00"),u'(x"1a"),u'(x"df"),u'(x"16"),u'(x"08"),u'(x"87"),u'(x"c1"),u'(x"ff"),u'(x"08"),u'(x"c1"),u'(x"c1"),u'(x"00"),u'(x"c1"),u'(x"01"),
u'(x"c9"),u'(x"01"),u'(x"0a"),u'(x"c1"),u'(x"00"),u'(x"c1"),u'(x"c1"),u'(x"00"),u'(x"c1"),u'(x"01"),u'(x"c9"),u'(x"01"),u'(x"00"),u'(x"87"),u'(x"c1"),u'(x"ff"),
u'(x"08"),u'(x"c1"),u'(x"c1"),u'(x"00"),u'(x"c1"),u'(x"01"),u'(x"c9"),u'(x"08"),u'(x"0a"),u'(x"c1"),u'(x"00"),u'(x"c1"),u'(x"c1"),u'(x"00"),u'(x"c1"),u'(x"01"),
u'(x"c9"),u'(x"08"),u'(x"00"),u'(x"87"),u'(x"87"),u'(x"77"),u'(x"b4"),u'(x"5f"),u'(x"08"),u'(x"87"),u'(x"c1"),u'(x"01"),u'(x"04"),u'(x"df"),u'(x"20"),u'(x"02"),
u'(x"03"),u'(x"df"),u'(x"20"),u'(x"02"),u'(x"c1"),u'(x"02"),u'(x"04"),u'(x"df"),u'(x"40"),u'(x"02"),u'(x"03"),u'(x"df"),u'(x"40"),u'(x"02"),u'(x"c1"),u'(x"04"),
u'(x"04"),u'(x"df"),u'(x"00"),u'(x"02"),u'(x"03"),u'(x"df"),u'(x"00"),u'(x"02"),u'(x"c1"),u'(x"08"),u'(x"04"),u'(x"df"),u'(x"00"),u'(x"02"),u'(x"03"),u'(x"df"),
u'(x"00"),u'(x"02"),u'(x"c1"),u'(x"10"),u'(x"02"),u'(x"f7"),u'(x"42"),u'(x"f7"),u'(x"4e"),u'(x"0a"),u'(x"c1"),u'(x"20"),u'(x"04"),u'(x"df"),u'(x"00"),u'(x"02"),
u'(x"03"),u'(x"df"),u'(x"00"),u'(x"02"),u'(x"87"),u'(x"c0"),u'(x"34"),u'(x"c0"),u'(x"c0"),u'(x"00"),u'(x"c0"),u'(x"00"),u'(x"48"),u'(x"b7"),u'(x"24"),u'(x"f7"),
u'(x"00"),u'(x"1e"),u'(x"df"),u'(x"1a"),u'(x"08"),u'(x"87"),u'(x"c1"),u'(x"ff"),u'(x"08"),u'(x"c1"),u'(x"c1"),u'(x"00"),u'(x"c1"),u'(x"01"),u'(x"c9"),u'(x"02"),
u'(x"0a"),u'(x"c1"),u'(x"00"),u'(x"c1"),u'(x"c1"),u'(x"00"),u'(x"c1"),u'(x"01"),u'(x"c9"),u'(x"02"),u'(x"00"),u'(x"87"),u'(x"c1"),u'(x"ff"),u'(x"08"),u'(x"c1"),
u'(x"c1"),u'(x"00"),u'(x"c1"),u'(x"01"),u'(x"c9"),u'(x"04"),u'(x"0a"),u'(x"c1"),u'(x"00"),u'(x"c1"),u'(x"c1"),u'(x"00"),u'(x"c1"),u'(x"01"),u'(x"c9"),u'(x"04"),
u'(x"00"),u'(x"87"),u'(x"c1"),u'(x"00"),u'(x"c1"),u'(x"e0"),u'(x"c1"),u'(x"c0"),u'(x"c1"),u'(x"40"),u'(x"c2"),u'(x"c8"),u'(x"87"),u'(x"f7"),u'(x"b8"),u'(x"c0"),
u'(x"44"),u'(x"f7"),u'(x"44"),u'(x"87"),u'(x"f7"),u'(x"aa"),u'(x"c0"),u'(x"42"),u'(x"f7"),u'(x"36"),u'(x"87"),u'(x"f7"),u'(x"9c"),u'(x"c0"),u'(x"43"),u'(x"f7"),
u'(x"28"),u'(x"87"),u'(x"f7"),u'(x"8e"),u'(x"c0"),u'(x"41"),u'(x"f7"),u'(x"1a"),u'(x"87"),u'(x"c1"),u'(x"14"),u'(x"f7"),u'(x"7c"),u'(x"c0"),u'(x"42"),u'(x"f7"),
u'(x"08"),u'(x"c1"),u'(x"f8"),u'(x"87"),u'(x"c1"),u'(x"14"),u'(x"f7"),u'(x"66"),u'(x"c0"),u'(x"41"),u'(x"f7"),u'(x"f2"),u'(x"c1"),u'(x"f8"),u'(x"87"),u'(x"c0"),
u'(x"0d"),u'(x"f7"),u'(x"e4"),u'(x"f7"),u'(x"3a"),u'(x"04"),u'(x"c0"),u'(x"0a"),u'(x"f7"),u'(x"d6"),u'(x"87"),u'(x"c0"),u'(x"1b"),u'(x"f7"),u'(x"cc"),u'(x"f7"),
u'(x"17"),u'(x"04"),u'(x"c0"),u'(x"4f"),u'(x"f7"),u'(x"be"),u'(x"c0"),u'(x"50"),u'(x"f7"),u'(x"b6"),u'(x"87"),u'(x"c0"),u'(x"1b"),u'(x"f7"),u'(x"ac"),u'(x"f7"),
u'(x"f7"),u'(x"04"),u'(x"c0"),u'(x"4f"),u'(x"f7"),u'(x"9e"),u'(x"c0"),u'(x"51"),u'(x"f7"),u'(x"96"),u'(x"87"),u'(x"c0"),u'(x"1b"),u'(x"f7"),u'(x"8c"),u'(x"f7"),
u'(x"d7"),u'(x"04"),u'(x"c0"),u'(x"4f"),u'(x"f7"),u'(x"7e"),u'(x"c0"),u'(x"52"),u'(x"f7"),u'(x"76"),u'(x"87"),u'(x"c0"),u'(x"1b"),u'(x"f7"),u'(x"6c"),u'(x"f7"),
u'(x"b7"),u'(x"04"),u'(x"c0"),u'(x"4f"),u'(x"f7"),u'(x"5e"),u'(x"c0"),u'(x"53"),u'(x"f7"),u'(x"56"),u'(x"87"),u'(x"f7"),u'(x"ae"),u'(x"05"),u'(x"c0"),u'(x"2b"),
u'(x"f7"),u'(x"46"),u'(x"87"),u'(x"87"),u'(x"f7"),u'(x"9c"),u'(x"03"),u'(x"f7"),u'(x"4c"),u'(x"87"),u'(x"f7"),u'(x"c8"),u'(x"c0"),u'(x"4d"),u'(x"f7"),u'(x"2a"),
u'(x"87"),u'(x"f7"),u'(x"82"),u'(x"05"),u'(x"c0"),u'(x"2e"),u'(x"f7"),u'(x"1a"),u'(x"87"),u'(x"f7"),u'(x"aa"),u'(x"c0"),u'(x"6e"),u'(x"f7"),u'(x"0c"),u'(x"87"),
u'(x"f7"),u'(x"64"),u'(x"05"),u'(x"c0"),u'(x"30"),u'(x"f7"),u'(x"fc"),u'(x"87"),u'(x"f7"),u'(x"8c"),u'(x"c0"),u'(x"70"),u'(x"f7"),u'(x"ee"),u'(x"87"),u'(x"f7"),
u'(x"46"),u'(x"05"),u'(x"c0"),u'(x"31"),u'(x"f7"),u'(x"de"),u'(x"87"),u'(x"f7"),u'(x"6e"),u'(x"c0"),u'(x"71"),u'(x"f7"),u'(x"d0"),u'(x"87"),u'(x"f7"),u'(x"28"),
u'(x"05"),u'(x"c0"),u'(x"32"),u'(x"f7"),u'(x"c0"),u'(x"87"),u'(x"f7"),u'(x"50"),u'(x"c0"),u'(x"72"),u'(x"f7"),u'(x"b2"),u'(x"87"),u'(x"f7"),u'(x"0a"),u'(x"05"),
u'(x"c0"),u'(x"33"),u'(x"f7"),u'(x"a2"),u'(x"87"),u'(x"f7"),u'(x"32"),u'(x"c0"),u'(x"73"),u'(x"f7"),u'(x"94"),u'(x"87"),u'(x"f7"),u'(x"ec"),u'(x"05"),u'(x"c0"),
u'(x"34"),u'(x"f7"),u'(x"84"),u'(x"87"),u'(x"f7"),u'(x"14"),u'(x"c0"),u'(x"74"),u'(x"f7"),u'(x"76"),u'(x"87"),u'(x"f7"),u'(x"ce"),u'(x"05"),u'(x"c0"),u'(x"35"),
u'(x"f7"),u'(x"66"),u'(x"87"),u'(x"f7"),u'(x"f6"),u'(x"c0"),u'(x"75"),u'(x"f7"),u'(x"58"),u'(x"87"),u'(x"f7"),u'(x"b0"),u'(x"05"),u'(x"c0"),u'(x"36"),u'(x"f7"),
u'(x"48"),u'(x"87"),u'(x"f7"),u'(x"d8"),u'(x"c0"),u'(x"76"),u'(x"f7"),u'(x"3a"),u'(x"87"),u'(x"f7"),u'(x"92"),u'(x"05"),u'(x"c0"),u'(x"37"),u'(x"f7"),u'(x"2a"),
u'(x"87"),u'(x"f7"),u'(x"ba"),u'(x"c0"),u'(x"77"),u'(x"f7"),u'(x"1c"),u'(x"87"),u'(x"f7"),u'(x"74"),u'(x"05"),u'(x"c0"),u'(x"38"),u'(x"f7"),u'(x"0c"),u'(x"87"),
u'(x"f7"),u'(x"9c"),u'(x"c0"),u'(x"78"),u'(x"f7"),u'(x"fe"),u'(x"87"),u'(x"f7"),u'(x"56"),u'(x"05"),u'(x"c0"),u'(x"39"),u'(x"f7"),u'(x"ee"),u'(x"87"),u'(x"f7"),
u'(x"7e"),u'(x"c0"),u'(x"79"),u'(x"f7"),u'(x"e0"),u'(x"87"),u'(x"87"),u'(x"87"),u'(x"c0"),u'(x"7f"),u'(x"f7"),u'(x"d2"),u'(x"87"),u'(x"87"),u'(x"f7"),u'(x"60"),
u'(x"c0"),u'(x"50"),u'(x"f7"),u'(x"c2"),u'(x"87"),u'(x"f7"),u'(x"52"),u'(x"c0"),u'(x"51"),u'(x"f7"),u'(x"b4"),u'(x"87"),u'(x"f7"),u'(x"44"),u'(x"c0"),u'(x"52"),
u'(x"f7"),u'(x"a6"),u'(x"87"),u'(x"f7"),u'(x"36"),u'(x"c0"),u'(x"53"),u'(x"f7"),u'(x"98"),u'(x"87"),u'(x"87"),u'(x"c0"),u'(x"1b"),u'(x"f7"),u'(x"8c"),u'(x"f7"),
u'(x"d7"),u'(x"0d"),u'(x"f7"),u'(x"df"),u'(x"05"),u'(x"c0"),u'(x"5b"),u'(x"f7"),u'(x"78"),u'(x"05"),u'(x"c0"),u'(x"4f"),u'(x"f7"),u'(x"6e"),u'(x"00"),u'(x"87"),
u'(x"c0"),u'(x"1b"),u'(x"f7"),u'(x"62"),u'(x"f7"),u'(x"ad"),u'(x"05"),u'(x"c0"),u'(x"4f"),u'(x"f7"),u'(x"54"),u'(x"87"),u'(x"c0"),u'(x"3f"),u'(x"f7"),u'(x"4a"),
u'(x"87"),u'(x"66"),u'(x"ba"),u'(x"c8"),u'(x"d6"),u'(x"e4"),u'(x"f2"),u'(x"08"),u'(x"1e"),u'(x"56"),u'(x"36"),u'(x"c8"),u'(x"76"),u'(x"96"),u'(x"b6"),u'(x"e2"),
u'(x"00"),u'(x"1e"),u'(x"3c"),u'(x"5a"),u'(x"78"),u'(x"96"),u'(x"b4"),u'(x"d2"),u'(x"f0"),u'(x"0e"),u'(x"2c"),u'(x"2e"),u'(x"30"),u'(x"3a"),u'(x"3c"),u'(x"4a"),
u'(x"58"),u'(x"f7"),u'(x"84"),u'(x"c0"),u'(x"00"),u'(x"c1"),u'(x"00"),u'(x"d0"),u'(x"45"),u'(x"01"),u'(x"fc"),u'(x"87"),u'(x"c0"),u'(x"d0"),u'(x"c0"),u'(x"f0"),
u'(x"05"),u'(x"20"),u'(x"f7"),u'(x"32"),u'(x"87"),u'(x"c0"),u'(x"be"),u'(x"c0"),u'(x"f0"),u'(x"07"),u'(x"20"),u'(x"f7"),u'(x"20"),u'(x"87"),u'(x"c0"),u'(x"ac"),
u'(x"c0"),u'(x"f0"),u'(x"04"),u'(x"20"),u'(x"f7"),u'(x"0e"),u'(x"87"),u'(x"c0"),u'(x"9a"),u'(x"c0"),u'(x"30"),u'(x"20"),u'(x"87"),u'(x"d7"),u'(x"92"),u'(x"28"),
u'(x"03"),u'(x"f7"),u'(x"28"),u'(x"88"),u'(x"c0"),u'(x"80"),u'(x"01"),u'(x"c0"),u'(x"c0"),u'(x"00"),u'(x"6e"),u'(x"c0"),u'(x"50"),u'(x"c1"),u'(x"41"),u'(x"6e"),
u'(x"d0"),u'(x"20"),u'(x"01"),u'(x"fc"),u'(x"87"),u'(x"66"),u'(x"26"),u'(x"c0"),u'(x"20"),u'(x"c1"),u'(x"38"),u'(x"10"),u'(x"01"),u'(x"fd"),u'(x"80"),u'(x"81"),
u'(x"87"),u'(x"66"),u'(x"26"),u'(x"c0"),u'(x"20"),u'(x"c0"),u'(x"3e"),u'(x"c0"),u'(x"c1"),u'(x"38"),u'(x"10"),u'(x"01"),u'(x"fd"),u'(x"80"),u'(x"81"),u'(x"87"),
u'(x"66"),u'(x"26"),u'(x"c0"),u'(x"20"),u'(x"01"),u'(x"c1"),u'(x"1e"),u'(x"10"),u'(x"01"),u'(x"fd"),u'(x"80"),u'(x"81"),u'(x"87"),u'(x"66"),u'(x"26"),u'(x"c0"),
u'(x"00"),u'(x"c1"),u'(x"00"),u'(x"d0"),u'(x"20"),u'(x"01"),u'(x"fc"),u'(x"f7"),u'(x"01"),u'(x"f8"),u'(x"f7"),u'(x"01"),u'(x"f6"),u'(x"37"),u'(x"f6"),u'(x"f7"),
u'(x"88"),u'(x"80"),u'(x"81"),u'(x"87"),u'(x"df"),u'(x"69"),u'(x"0a"),u'(x"03"),u'(x"f7"),u'(x"01"),u'(x"45"),u'(x"87"),u'(x"37"),u'(x"3f"),u'(x"87"),u'(x"f7"),
u'(x"ca"),u'(x"ca"),u'(x"f7"),u'(x"c8"),u'(x"c8"),u'(x"f7"),u'(x"c6"),u'(x"c5"),u'(x"f7"),u'(x"c6"),u'(x"c5"),u'(x"f7"),u'(x"bc"),u'(x"bb"),u'(x"87"),u'(x"f7"),
u'(x"ac"),u'(x"a8"),u'(x"f7"),u'(x"aa"),u'(x"a6"),u'(x"f7"),u'(x"a7"),u'(x"a4"),u'(x"f7"),u'(x"a7"),u'(x"a4"),u'(x"f7"),u'(x"9d"),u'(x"9a"),u'(x"f7"),u'(x"ca"),
u'(x"87"),u'(x"37"),u'(x"f3"),u'(x"87"),u'(x"f7"),u'(x"01"),u'(x"fa"),u'(x"87"),u'(x"37"),u'(x"f4"),u'(x"87"),u'(x"f7"),u'(x"72"),u'(x"f7"),u'(x"ac"),u'(x"87"),
u'(x"b7"),u'(x"68"),u'(x"f7"),u'(x"a2"),u'(x"87"),u'(x"b7"),u'(x"62"),u'(x"f7"),u'(x"98"),u'(x"87"),u'(x"f7"),u'(x"c1"),u'(x"0c"),u'(x"f7"),u'(x"62"),u'(x"4c"),
u'(x"03"),u'(x"b7"),u'(x"46"),u'(x"02"),u'(x"f7"),u'(x"ec"),u'(x"37"),u'(x"44"),u'(x"87"),u'(x"f7"),u'(x"3a"),u'(x"f7"),u'(x"70"),u'(x"87"),u'(x"f7"),u'(x"01"),
u'(x"2e"),u'(x"f7"),u'(x"3a"),u'(x"24"),u'(x"03"),u'(x"b7"),u'(x"1e"),u'(x"02"),u'(x"f7"),u'(x"c4"),u'(x"37"),u'(x"1c"),u'(x"87"),u'(x"87"),u'(x"87"),u'(x"f7"),
u'(x"77"),u'(x"07"),u'(x"c0"),u'(x"08"),u'(x"c0"),u'(x"f0"),u'(x"01"),u'(x"02"),u'(x"87"),u'(x"f7"),u'(x"01"),u'(x"f8"),u'(x"f7"),u'(x"01"),u'(x"ee"),u'(x"87"),
u'(x"f7"),u'(x"01"),u'(x"e6"),u'(x"03"),u'(x"f7"),u'(x"e0"),u'(x"02"),u'(x"f7"),u'(x"e0"),u'(x"37"),u'(x"de"),u'(x"87"),u'(x"f7"),u'(x"0e"),u'(x"c1"),u'(x"00"),
u'(x"d0"),u'(x"20"),u'(x"01"),u'(x"fc"),u'(x"87"),u'(x"f7"),u'(x"fc"),u'(x"c1"),u'(x"ba"),u'(x"c1"),u'(x"41"),u'(x"6e"),u'(x"d0"),u'(x"20"),u'(x"01"),u'(x"fc"),
u'(x"87"),u'(x"f7"),u'(x"24"),u'(x"07"),u'(x"f7"),u'(x"b0"),u'(x"9e"),u'(x"0a"),u'(x"f7"),u'(x"98"),u'(x"09"),u'(x"f7"),u'(x"01"),u'(x"90"),u'(x"03"),u'(x"f7"),
u'(x"8a"),u'(x"02"),u'(x"f7"),u'(x"8a"),u'(x"37"),u'(x"88"),u'(x"87"),u'(x"f7"),u'(x"e7"),u'(x"03"),u'(x"f7"),u'(x"76"),u'(x"87"),u'(x"c0"),u'(x"1b"),u'(x"f7"),
u'(x"88"),u'(x"c0"),u'(x"2f"),u'(x"f7"),u'(x"80"),u'(x"c0"),u'(x"5a"),u'(x"f7"),u'(x"78"),u'(x"87"),u'(x"77"),u'(x"68"),u'(x"a6"),u'(x"f7"),u'(x"8c"),u'(x"02"),
u'(x"c0"),u'(x"48"),u'(x"c0"),u'(x"00"),u'(x"6e"),u'(x"01"),u'(x"c1"),u'(x"c1"),u'(x"42"),u'(x"0c"),u'(x"60"),u'(x"42"),u'(x"fd"),u'(x"ca"),u'(x"20"),u'(x"f7"),
u'(x"01"),u'(x"bc"),u'(x"03"),u'(x"f7"),u'(x"b6"),u'(x"ea"),u'(x"82"),u'(x"87"),u'(x"f7"),u'(x"ac"),u'(x"16"),u'(x"f7"),u'(x"50"),u'(x"37"),u'(x"16"),u'(x"87"),
u'(x"f7"),u'(x"9c"),u'(x"06"),u'(x"f7"),u'(x"40"),u'(x"37"),u'(x"06"),u'(x"87"),u'(x"f7"),u'(x"8c"),u'(x"fa"),u'(x"f7"),u'(x"30"),u'(x"37"),u'(x"f6"),u'(x"87"),
u'(x"f7"),u'(x"7c"),u'(x"ea"),u'(x"f7"),u'(x"20"),u'(x"37"),u'(x"e6"),u'(x"87"),u'(x"f7"),u'(x"6c"),u'(x"d6"),u'(x"f7"),u'(x"68"),u'(x"d4"),u'(x"f7"),u'(x"0a"),
u'(x"37"),u'(x"d0"),u'(x"87"),u'(x"f7"),u'(x"00"),u'(x"f7"),u'(x"40"),u'(x"05"),u'(x"f7"),u'(x"6e"),u'(x"c1"),u'(x"00"),u'(x"1b"),u'(x"f7"),u'(x"01"),u'(x"2e"),
u'(x"07"),u'(x"f7"),u'(x"7a"),u'(x"01"),u'(x"81"),u'(x"c0"),u'(x"00"),u'(x"10"),u'(x"f7"),u'(x"02"),u'(x"18"),u'(x"05"),u'(x"f7"),u'(x"03"),u'(x"10"),u'(x"01"),
u'(x"07"),u'(x"f7"),u'(x"24"),u'(x"c0"),u'(x"00"),u'(x"c1"),u'(x"00"),u'(x"00"),u'(x"d0"),u'(x"20"),u'(x"01"),u'(x"fc"),u'(x"00"),u'(x"37"),u'(x"76"),u'(x"87"),
u'(x"f7"),u'(x"a6"),u'(x"f7"),u'(x"e6"),u'(x"06"),u'(x"c1"),u'(x"5e"),u'(x"c1"),u'(x"41"),u'(x"6e"),u'(x"1d"),u'(x"f7"),u'(x"01"),u'(x"d2"),u'(x"09"),u'(x"01"),
u'(x"81"),u'(x"c0"),u'(x"46"),u'(x"c0"),u'(x"c0"),u'(x"00"),u'(x"6e"),u'(x"10"),u'(x"f7"),u'(x"02"),u'(x"b8"),u'(x"11"),u'(x"c0"),u'(x"30"),u'(x"c0"),u'(x"c0"),
u'(x"00"),u'(x"6e"),u'(x"c1"),u'(x"24"),u'(x"c1"),u'(x"41"),u'(x"6e"),u'(x"00"),u'(x"d0"),u'(x"20"),u'(x"01"),u'(x"fc"),u'(x"00"),u'(x"37"),u'(x"16"),u'(x"87"),
u'(x"a6"),u'(x"f7"),u'(x"06"),u'(x"18"),u'(x"23"),u'(x"c0"),u'(x"10"),u'(x"c0"),u'(x"00"),u'(x"6e"),u'(x"c1"),u'(x"06"),u'(x"c1"),u'(x"84"),u'(x"c1"),u'(x"41"),
u'(x"6e"),u'(x"c2"),u'(x"f6"),u'(x"c2"),u'(x"c2"),u'(x"e0"),u'(x"c2"),u'(x"c2"),u'(x"82"),u'(x"6e"),u'(x"42"),u'(x"03"),u'(x"60"),u'(x"42"),u'(x"fd"),u'(x"c0"),
u'(x"c0"),u'(x"c8"),u'(x"20"),u'(x"02"),u'(x"fa"),u'(x"f7"),u'(x"01"),u'(x"c0"),u'(x"82"),u'(x"87"),u'(x"a6"),u'(x"f7"),u'(x"b2"),u'(x"c4"),u'(x"26"),u'(x"c0"),
u'(x"ba"),u'(x"c0"),u'(x"a6"),u'(x"c0"),u'(x"c0"),u'(x"01"),u'(x"c1"),u'(x"30"),u'(x"c2"),u'(x"ac"),u'(x"c2"),u'(x"94"),u'(x"81"),u'(x"01"),u'(x"81"),u'(x"c1"),
u'(x"c0"),u'(x"41"),u'(x"6e"),u'(x"00"),u'(x"6e"),u'(x"c2"),u'(x"90"),u'(x"c2"),u'(x"82"),u'(x"6e"),u'(x"50"),u'(x"42"),u'(x"fd"),u'(x"d0"),u'(x"20"),u'(x"80"),
u'(x"02"),u'(x"fb"),u'(x"f7"),u'(x"01"),u'(x"66"),u'(x"82"),u'(x"87"),u'(x"a6"),u'(x"c2"),u'(x"58"),u'(x"c2"),u'(x"82"),u'(x"6e"),u'(x"f7"),u'(x"8c"),u'(x"01"),
u'(x"c1"),u'(x"dc"),u'(x"c1"),u'(x"d8"),u'(x"42"),u'(x"02"),u'(x"81"),u'(x"03"),u'(x"50"),u'(x"42"),u'(x"fd"),u'(x"d0"),u'(x"20"),u'(x"02"),u'(x"fc"),u'(x"82"),
u'(x"87"),u'(x"a6"),u'(x"c2"),u'(x"24"),u'(x"c2"),u'(x"82"),u'(x"6e"),u'(x"f7"),u'(x"58"),u'(x"01"),u'(x"c1"),u'(x"a8"),u'(x"c1"),u'(x"a4"),u'(x"42"),u'(x"01"),
u'(x"81"),u'(x"d0"),u'(x"20"),u'(x"01"),u'(x"fc"),u'(x"82"),u'(x"87"),u'(x"c1"),u'(x"00"),u'(x"40"),u'(x"f7"),u'(x"12"),u'(x"57"),u'(x"07"),u'(x"fa"),u'(x"87"),
u'(x"1b"),u'(x"3f"),u'(x"3b"),u'(x"63"),u'(x"f7"),u'(x"04"),u'(x"87"),u'(x"f7"),u'(x"00"),u'(x"5a"),u'(x"06"),u'(x"c0"),u'(x"d6"),u'(x"c0"),u'(x"30"),u'(x"02"),
u'(x"0c"),u'(x"f7"),u'(x"03"),u'(x"46"),u'(x"08"),u'(x"c0"),u'(x"50"),u'(x"c0"),u'(x"30"),u'(x"02"),u'(x"c0"),u'(x"c0"),u'(x"fb"),u'(x"87"),u'(x"00"),u'(x"37"),
u'(x"2a"),u'(x"3a"),u'(x"01"),u'(x"6e"),u'(x"c1"),u'(x"14"),u'(x"04"),u'(x"f7"),u'(x"01"),u'(x"10"),u'(x"2e"),u'(x"c1"),u'(x"01"),u'(x"04"),u'(x"f7"),u'(x"01"),
u'(x"05"),u'(x"27"),u'(x"c1"),u'(x"03"),u'(x"06"),u'(x"f7"),u'(x"01"),u'(x"f9"),u'(x"f7"),u'(x"66"),u'(x"1e"),u'(x"c1"),u'(x"04"),u'(x"04"),u'(x"f7"),u'(x"01"),
u'(x"e3"),u'(x"17"),u'(x"c1"),u'(x"06"),u'(x"06"),u'(x"f7"),u'(x"01"),u'(x"da"),u'(x"37"),u'(x"60"),u'(x"0e"),u'(x"c1"),u'(x"07"),u'(x"04"),u'(x"f7"),u'(x"01"),
u'(x"c4"),u'(x"07"),u'(x"c1"),u'(x"19"),u'(x"04"),u'(x"df"),u'(x"80"),u'(x"02"),u'(x"00"),u'(x"80"),u'(x"80"),u'(x"c3"),u'(x"87"),u'(x"00"),u'(x"37"),u'(x"ac"),
u'(x"41"),u'(x"01"),u'(x"6e"),u'(x"c1"),u'(x"02"),u'(x"04"),u'(x"f7"),u'(x"01"),u'(x"87"),u'(x"35"),u'(x"c1"),u'(x"14"),u'(x"04"),u'(x"f7"),u'(x"00"),u'(x"84"),
u'(x"2e"),u'(x"c1"),u'(x"01"),u'(x"04"),u'(x"f7"),u'(x"00"),u'(x"79"),u'(x"27"),u'(x"c1"),u'(x"03"),u'(x"06"),u'(x"f7"),u'(x"00"),u'(x"6d"),u'(x"f7"),u'(x"da"),
u'(x"1e"),u'(x"c1"),u'(x"04"),u'(x"04"),u'(x"f7"),u'(x"00"),u'(x"57"),u'(x"17"),u'(x"c1"),u'(x"06"),u'(x"06"),u'(x"f7"),u'(x"00"),u'(x"4e"),u'(x"37"),u'(x"d4"),
u'(x"0e"),u'(x"c1"),u'(x"07"),u'(x"04"),u'(x"f7"),u'(x"00"),u'(x"38"),u'(x"07"),u'(x"c1"),u'(x"19"),u'(x"04"),u'(x"df"),u'(x"80"),u'(x"02"),u'(x"00"),u'(x"80"),
u'(x"80"),u'(x"bc"),u'(x"87"),u'(x"00"),u'(x"37"),u'(x"20"),u'(x"43"),u'(x"01"),u'(x"6e"),u'(x"c1"),u'(x"00"),u'(x"03"),u'(x"37"),u'(x"9a"),u'(x"38"),u'(x"c1"),
u'(x"01"),u'(x"04"),u'(x"f7"),u'(x"01"),u'(x"8c"),u'(x"31"),u'(x"c1"),u'(x"04"),u'(x"04"),u'(x"f7"),u'(x"02"),u'(x"7e"),u'(x"2a"),u'(x"c1"),u'(x"05"),u'(x"04"),
u'(x"f7"),u'(x"04"),u'(x"70"),u'(x"23"),u'(x"c1"),u'(x"07"),u'(x"04"),u'(x"f7"),u'(x"08"),u'(x"62"),u'(x"1c"),u'(x"c1"),u'(x"16"),u'(x"04"),u'(x"f7"),u'(x"01"),
u'(x"54"),u'(x"15"),u'(x"c1"),u'(x"18"),u'(x"04"),u'(x"f7"),u'(x"02"),u'(x"46"),u'(x"0e"),u'(x"c1"),u'(x"19"),u'(x"04"),u'(x"f7"),u'(x"04"),u'(x"38"),u'(x"07"),
u'(x"c1"),u'(x"1b"),u'(x"04"),u'(x"f7"),u'(x"08"),u'(x"2a"),u'(x"00"),u'(x"80"),u'(x"80"),u'(x"ba"),u'(x"87"),u'(x"f7"),u'(x"05"),u'(x"92"),u'(x"05"),u'(x"f7"),
u'(x"06"),u'(x"8a"),u'(x"12"),u'(x"47"),u'(x"c0"),u'(x"1b"),u'(x"f7"),u'(x"1a"),u'(x"c0"),u'(x"5b"),u'(x"f7"),u'(x"12"),u'(x"c0"),u'(x"30"),u'(x"f7"),u'(x"0a"),
u'(x"c0"),u'(x"6e"),u'(x"f7"),u'(x"02"),u'(x"36"),u'(x"c0"),u'(x"1b"),u'(x"f7"),u'(x"f8"),u'(x"c0"),u'(x"5b"),u'(x"f7"),u'(x"f0"),u'(x"c1"),u'(x"ce"),u'(x"00"),
u'(x"c0"),u'(x"80"),u'(x"c1"),u'(x"0a"),u'(x"fc"),u'(x"c1"),u'(x"3a"),u'(x"c0"),u'(x"04"),u'(x"c0"),u'(x"30"),u'(x"f7"),u'(x"d0"),u'(x"40"),u'(x"f7"),u'(x"ca"),
u'(x"c0"),u'(x"3b"),u'(x"f7"),u'(x"c2"),u'(x"c1"),u'(x"a4"),u'(x"00"),u'(x"c0"),u'(x"80"),u'(x"c1"),u'(x"0a"),u'(x"fc"),u'(x"c1"),u'(x"3a"),u'(x"c0"),u'(x"04"),
u'(x"c0"),u'(x"30"),u'(x"f7"),u'(x"a2"),u'(x"40"),u'(x"f7"),u'(x"9c"),u'(x"c0"),u'(x"52"),u'(x"f7"),u'(x"94"),u'(x"87"),u'(x"c0"),u'(x"f2"),u'(x"c0"),u'(x"0f"),
u'(x"c1"),u'(x"ec"),u'(x"c1"),u'(x"0b"),u'(x"01"),u'(x"09"),u'(x"37"),u'(x"6c"),u'(x"77"),u'(x"6a"),u'(x"01"),u'(x"81"),u'(x"77"),u'(x"64"),u'(x"09"),u'(x"f7"),
u'(x"01"),u'(x"58"),u'(x"f7"),u'(x"18"),u'(x"54"),u'(x"f7"),u'(x"18"),u'(x"50"),u'(x"c0"),u'(x"01"),u'(x"37"),u'(x"34"),u'(x"37"),u'(x"34"),u'(x"f7"),u'(x"6a"),
u'(x"37"),u'(x"30"),u'(x"87"),u'(x"f7"),u'(x"00"),u'(x"a2"),u'(x"09"),u'(x"c1"),u'(x"10"),u'(x"40"),u'(x"f7"),u'(x"32"),u'(x"57"),u'(x"24"),u'(x"fa"),u'(x"0d"),
u'(x"f7"),u'(x"01"),u'(x"88"),u'(x"09"),u'(x"c1"),u'(x"fc"),u'(x"40"),u'(x"f7"),u'(x"18"),u'(x"57"),u'(x"10"),u'(x"fa"),u'(x"00"),u'(x"87"),u'(x"1b"),u'(x"33"),
u'(x"31"),u'(x"31"),u'(x"31"),u'(x"32"),u'(x"31"),u'(x"32"),u'(x"31"),u'(x"30"),u'(x"1b"),u'(x"32"),u'(x"31"),u'(x"31"),u'(x"31"),u'(x"32"),u'(x"31"),u'(x"32"),
u'(x"31"),u'(x"30"),u'(x"77"),u'(x"d8"),u'(x"87"),u'(x"66"),u'(x"d7"),u'(x"c0"),u'(x"01"),u'(x"03"),u'(x"f7"),u'(x"01"),u'(x"b6"),u'(x"d7"),u'(x"b2"),u'(x"50"),
u'(x"03"),u'(x"f7"),u'(x"50"),u'(x"a8"),u'(x"c0"),u'(x"a0"),u'(x"17"),u'(x"01"),u'(x"04"),u'(x"f7"),u'(x"01"),u'(x"94"),u'(x"f7"),u'(x"17"),u'(x"18"),u'(x"04"),
u'(x"f7"),u'(x"18"),u'(x"86"),u'(x"f0"),u'(x"f7"),u'(x"fe"),u'(x"0a"),u'(x"37"),u'(x"8e"),u'(x"04"),u'(x"c0"),u'(x"88"),u'(x"37"),u'(x"70"),u'(x"c0"),u'(x"7c"),
u'(x"c0"),u'(x"c0"),u'(x"c0"),u'(x"00"),u'(x"6e"),u'(x"c1"),u'(x"62"),u'(x"c1"),u'(x"c1"),u'(x"40"),u'(x"81"),u'(x"87"),u'(x"a6"),u'(x"66"),u'(x"26"),u'(x"c1"),
u'(x"5a"),u'(x"40"),u'(x"c0"),u'(x"c1"),u'(x"c0"),u'(x"41"),u'(x"6e"),u'(x"00"),u'(x"6e"),u'(x"c2"),u'(x"48"),u'(x"c2"),u'(x"82"),u'(x"6e"),u'(x"50"),u'(x"42"),
u'(x"fd"),u'(x"d0"),u'(x"20"),u'(x"02"),u'(x"fc"),u'(x"c1"),u'(x"2e"),u'(x"40"),u'(x"c0"),u'(x"c1"),u'(x"20"),u'(x"c0"),u'(x"20"),u'(x"c2"),u'(x"20"),u'(x"c2"),
u'(x"20"),u'(x"50"),u'(x"42"),u'(x"fd"),u'(x"08"),u'(x"80"),u'(x"81"),u'(x"82"),u'(x"87"),u'(x"a6"),u'(x"66"),u'(x"26"),u'(x"c1"),u'(x"02"),u'(x"40"),u'(x"c1"),
u'(x"c1"),u'(x"c0"),u'(x"41"),u'(x"6e"),u'(x"00"),u'(x"6e"),u'(x"c2"),u'(x"ec"),u'(x"c2"),u'(x"c2"),u'(x"82"),u'(x"6e"),u'(x"60"),u'(x"42"),u'(x"fd"),u'(x"e0"),
u'(x"20"),u'(x"02"),u'(x"fc"),u'(x"c1"),u'(x"d4"),u'(x"40"),u'(x"c1"),u'(x"c1"),u'(x"20"),u'(x"c0"),u'(x"20"),u'(x"c2"),u'(x"c2"),u'(x"c2"),u'(x"c2"),u'(x"20"),
u'(x"60"),u'(x"42"),u'(x"fd"),u'(x"20"),u'(x"80"),u'(x"81"),u'(x"82"),u'(x"87"),u'(x"f7"),u'(x"a0"),u'(x"17"),u'(x"f7"),u'(x"ff"),u'(x"14"),u'(x"d7"),u'(x"90"),
u'(x"50"),u'(x"10"),u'(x"f7"),u'(x"84"),u'(x"94"),u'(x"07"),u'(x"f7"),u'(x"01"),u'(x"7e"),u'(x"f7"),u'(x"01"),u'(x"74"),u'(x"05"),u'(x"f7"),u'(x"1a"),u'(x"f7"),
u'(x"01"),u'(x"6c"),u'(x"37"),u'(x"6c"),u'(x"f7"),u'(x"9e"),u'(x"87"),u'(x"f7"),u'(x"be"),u'(x"d7"),u'(x"64"),u'(x"30"),u'(x"09"),u'(x"57"),u'(x"5f"),u'(x"06"),
u'(x"57"),u'(x"7f"),u'(x"03"),u'(x"c1"),u'(x"5f"),u'(x"0a"),u'(x"d7"),u'(x"4a"),u'(x"41"),u'(x"06"),u'(x"57"),u'(x"24"),u'(x"03"),u'(x"c1"),u'(x"1e"),u'(x"00"),
u'(x"f7"),u'(x"a1"),u'(x"14"),u'(x"26"),u'(x"66"),u'(x"a6"),u'(x"02"),u'(x"c0"),u'(x"1a"),u'(x"c0"),u'(x"00"),u'(x"6e"),u'(x"01"),u'(x"c1"),u'(x"c1"),u'(x"42"),
u'(x"03"),u'(x"60"),u'(x"42"),u'(x"fd"),u'(x"82"),u'(x"81"),u'(x"80"),u'(x"50"),u'(x"c8"),u'(x"02"),u'(x"c0"),u'(x"d7"),u'(x"f6"),u'(x"50"),u'(x"01"),u'(x"07"),
u'(x"f7"),u'(x"62"),u'(x"08"),u'(x"f7"),u'(x"01"),u'(x"e8"),u'(x"04"),u'(x"f7"),u'(x"01"),u'(x"dc"),u'(x"00"),u'(x"87"),u'(x"57"),u'(x"20"),u'(x"08"),u'(x"40"),
u'(x"c0"),u'(x"00"),u'(x"ae"),u'(x"c0"),u'(x"02"),u'(x"c8"),u'(x"01"),u'(x"87"),u'(x"87"),u'(x"87"),u'(x"df"),u'(x"69"),u'(x"0a"),u'(x"09"),u'(x"c1"),u'(x"60"),
u'(x"40"),u'(x"f7"),u'(x"c4"),u'(x"57"),u'(x"6e"),u'(x"fa"),u'(x"87"),u'(x"c1"),u'(x"6e"),u'(x"40"),u'(x"f7"),u'(x"b2"),u'(x"57"),u'(x"7c"),u'(x"fa"),u'(x"87"),
u'(x"76"),u'(x"31"),u'(x"30"),u'(x"70"),u'(x"70"),u'(x"30"),u'(x"31"),u'(x"76"),u'(x"31"),u'(x"35"),u'(x"70"),u'(x"70"),u'(x"30"),u'(x"31"),u'(x"f7"),u'(x"01"),
u'(x"6e"),u'(x"f7"),u'(x"a4"),u'(x"37"),u'(x"6a"),u'(x"87"),u'(x"c0"),u'(x"60"),u'(x"c1"),u'(x"02"),u'(x"01"),u'(x"c1"),u'(x"c0"),u'(x"50"),u'(x"c0"),u'(x"00"),
u'(x"20"),u'(x"c0"),u'(x"05"),u'(x"f7"),u'(x"28"),u'(x"44"),u'(x"0a"),u'(x"04"),u'(x"f7"),u'(x"50"),u'(x"3a"),u'(x"05"),u'(x"b7"),u'(x"34"),u'(x"81"),u'(x"c9"),
u'(x"f0"),u'(x"f7"),u'(x"64"),u'(x"37"),u'(x"2a"),u'(x"87"),u'(x"f7"),u'(x"94"),u'(x"03"),u'(x"f7"),u'(x"01"),u'(x"18"),u'(x"f7"),u'(x"8e"),u'(x"07"),u'(x"f7"),
u'(x"0a"),u'(x"1c"),u'(x"0f"),u'(x"f7"),u'(x"ae"),u'(x"10"),u'(x"f7"),u'(x"fc"),u'(x"0a"),u'(x"08"),u'(x"f7"),u'(x"f4"),u'(x"04"),u'(x"04"),u'(x"03"),u'(x"f7"),
u'(x"96"),u'(x"04"),u'(x"f7"),u'(x"01"),u'(x"e2"),u'(x"00"),u'(x"37"),u'(x"e4"),u'(x"87"),u'(x"f7"),u'(x"01"),u'(x"d8"),u'(x"f7"),u'(x"0e"),u'(x"37"),u'(x"d4"),
u'(x"87"),u'(x"f7"),u'(x"d3"),u'(x"d2"),u'(x"87"),u'(x"f7"),u'(x"ca"),u'(x"ca"),u'(x"87"),u'(x"f7"),u'(x"00"),u'(x"4c"),u'(x"37"),u'(x"b8"),u'(x"87"),u'(x"f7"),
u'(x"19"),u'(x"03"),u'(x"f7"),u'(x"5e"),u'(x"09"),u'(x"57"),u'(x"20"),u'(x"06"),u'(x"57"),u'(x"7f"),u'(x"03"),u'(x"f7"),u'(x"34"),u'(x"00"),u'(x"87"),u'(x"57"),
u'(x"40"),u'(x"20"),u'(x"57"),u'(x"7f"),u'(x"1d"),u'(x"c1"),u'(x"c0"),u'(x"c1"),u'(x"c1"),u'(x"ee"),u'(x"41"),u'(x"f7"),u'(x"f4"),u'(x"04"),u'(x"f7"),u'(x"00"),
u'(x"03"),u'(x"f7"),u'(x"01"),u'(x"f8"),u'(x"f7"),u'(x"e4"),u'(x"f4"),u'(x"f7"),u'(x"f0"),u'(x"03"),u'(x"f7"),u'(x"01"),u'(x"e8"),u'(x"c9"),u'(x"f7"),u'(x"00"),
u'(x"e2"),u'(x"26"),u'(x"57"),u'(x"30"),u'(x"19"),u'(x"57"),u'(x"39"),u'(x"16"),u'(x"c0"),u'(x"b8"),u'(x"17"),u'(x"0e"),u'(x"02"),u'(x"c0"),u'(x"0e"),u'(x"02"),
u'(x"6e"),u'(x"c2"),u'(x"c2"),u'(x"c2"),u'(x"02"),u'(x"6e"),u'(x"02"),u'(x"6e"),u'(x"c1"),u'(x"f0"),u'(x"42"),u'(x"b0"),u'(x"6e"),u'(x"0a"),u'(x"57"),u'(x"3b"),
u'(x"04"),u'(x"f7"),u'(x"02"),u'(x"84"),u'(x"03"),u'(x"57"),u'(x"3f"),u'(x"00"),u'(x"87"),u'(x"f7"),u'(x"00"),u'(x"8c"),u'(x"87"),u'(x"f7"),u'(x"00"),u'(x"84"),
u'(x"87"),u'(x"37"),u'(x"66"),u'(x"c0"),u'(x"6e"),u'(x"10"),u'(x"17"),u'(x"7e"),u'(x"fc"),u'(x"57"),u'(x"3a"),u'(x"04"),u'(x"f7"),u'(x"04"),u'(x"66"),u'(x"0c"),
u'(x"57"),u'(x"30"),u'(x"09"),u'(x"57"),u'(x"7e"),u'(x"06"),u'(x"f7"),u'(x"02"),u'(x"52"),u'(x"f7"),u'(x"28"),u'(x"00"),u'(x"87"),u'(x"d7"),u'(x"2d"),u'(x"23"),
u'(x"1e"),u'(x"57"),u'(x"38"),u'(x"03"),u'(x"f7"),u'(x"b6"),u'(x"46"),u'(x"57"),u'(x"33"),u'(x"03"),u'(x"f7"),u'(x"c0"),u'(x"40"),u'(x"57"),u'(x"34"),u'(x"03"),
u'(x"f7"),u'(x"c6"),u'(x"3a"),u'(x"57"),u'(x"35"),u'(x"03"),u'(x"f7"),u'(x"de"),u'(x"34"),u'(x"57"),u'(x"36"),u'(x"03"),u'(x"f7"),u'(x"c0"),u'(x"2e"),u'(x"d7"),
u'(x"e9"),u'(x"28"),u'(x"05"),u'(x"77"),u'(x"6e"),u'(x"77"),u'(x"6c"),u'(x"25"),u'(x"d7"),u'(x"d7"),u'(x"29"),u'(x"05"),u'(x"77"),u'(x"5d"),u'(x"77"),u'(x"5a"),
u'(x"1c"),u'(x"d7"),u'(x"c5"),u'(x"59"),u'(x"18"),u'(x"f7"),u'(x"ab"),u'(x"15"),u'(x"f7"),u'(x"a6"),u'(x"05"),u'(x"c1"),u'(x"1f"),u'(x"77"),u'(x"9c"),u'(x"10"),
u'(x"c1"),u'(x"1f"),u'(x"77"),u'(x"28"),u'(x"c1"),u'(x"8e"),u'(x"77"),u'(x"1c"),u'(x"37"),u'(x"86"),u'(x"f7"),u'(x"52"),u'(x"00"),u'(x"f7"),u'(x"00"),u'(x"a4"),
u'(x"87"),u'(x"57"),u'(x"1b"),u'(x"01"),u'(x"12"),u'(x"77"),u'(x"7d"),u'(x"40"),u'(x"c0"),u'(x"80"),u'(x"c0"),u'(x"00"),u'(x"ae"),u'(x"17"),u'(x"40"),u'(x"03"),
u'(x"37"),u'(x"80"),u'(x"04"),u'(x"c8"),u'(x"f7"),u'(x"00"),u'(x"76"),u'(x"87"),u'(x"f7"),u'(x"00"),u'(x"6e"),u'(x"87"),u'(x"f7"),u'(x"00"),u'(x"66"),u'(x"87"),
u'(x"f7"),u'(x"00"),u'(x"5e"),u'(x"87"),u'(x"f7"),u'(x"00"),u'(x"56"),u'(x"87"),u'(x"f7"),u'(x"00"),u'(x"4e"),u'(x"87"),u'(x"f7"),u'(x"00"),u'(x"46"),u'(x"87"),
u'(x"f7"),u'(x"00"),u'(x"3e"),u'(x"87"),u'(x"f7"),u'(x"00"),u'(x"36"),u'(x"87"),u'(x"a6"),u'(x"66"),u'(x"00"),u'(x"c1"),u'(x"00"),u'(x"c2"),u'(x"00"),u'(x"11"),
u'(x"81"),u'(x"fd"),u'(x"81"),u'(x"82"),u'(x"87"),u'(x"df"),u'(x"e0"),u'(x"fe"),u'(x"c0"),u'(x"72"),u'(x"c1"),u'(x"6c"),u'(x"01"),u'(x"02"),u'(x"00"),u'(x"1e"),
u'(x"f7"),u'(x"5c"),u'(x"80"),u'(x"17"),u'(x"80"),u'(x"01"),u'(x"00"),u'(x"37"),u'(x"54"),u'(x"c0"),u'(x"40"),u'(x"01"),u'(x"c1"),u'(x"00"),u'(x"f7"),u'(x"42"),
u'(x"0d"),u'(x"d7"),u'(x"3a"),u'(x"10"),u'(x"09"),u'(x"f7"),u'(x"35"),u'(x"06"),u'(x"c0"),u'(x"11"),u'(x"f7"),u'(x"52"),u'(x"37"),u'(x"26"),u'(x"df"),u'(x"00"),
u'(x"fe"),u'(x"87"),u'(x"df"),u'(x"e0"),u'(x"fe"),u'(x"c0"),u'(x"1c"),u'(x"c1"),u'(x"16"),u'(x"01"),u'(x"02"),u'(x"00"),u'(x"0c"),u'(x"80"),u'(x"17"),u'(x"20"),
u'(x"01"),u'(x"00"),u'(x"37"),u'(x"02"),u'(x"c0"),u'(x"c0"),u'(x"01"),u'(x"c1"),u'(x"00"),u'(x"df"),u'(x"00"),u'(x"fe"),u'(x"87"),u'(x"57"),u'(x"14"),u'(x"09"),
u'(x"f7"),u'(x"4f"),u'(x"03"),u'(x"37"),u'(x"4a"),u'(x"0d"),u'(x"37"),u'(x"45"),u'(x"0a"),u'(x"57"),u'(x"12"),u'(x"02"),u'(x"37"),u'(x"3a"),u'(x"57"),u'(x"59"),
u'(x"02"),u'(x"37"),u'(x"31"),u'(x"87"),u'(x"40"),u'(x"57"),u'(x"14"),u'(x"0d"),u'(x"f7"),u'(x"1f"),u'(x"05"),u'(x"f7"),u'(x"01"),u'(x"18"),u'(x"00"),u'(x"24"),
u'(x"f7"),u'(x"01"),u'(x"0f"),u'(x"00"),u'(x"1f"),u'(x"57"),u'(x"12"),u'(x"05"),u'(x"f7"),u'(x"01"),u'(x"00"),u'(x"00"),u'(x"17"),u'(x"57"),u'(x"59"),u'(x"05"),
u'(x"f7"),u'(x"01"),u'(x"f1"),u'(x"00"),u'(x"0f"),u'(x"57"),u'(x"58"),u'(x"0c"),u'(x"f7"),u'(x"e4"),u'(x"04"),u'(x"37"),u'(x"de"),u'(x"00"),u'(x"05"),u'(x"f7"),
u'(x"01"),u'(x"d4"),u'(x"00"),u'(x"00"),u'(x"87"),u'(x"f7"),u'(x"c4"),u'(x"08"),u'(x"f7"),u'(x"66"),u'(x"37"),u'(x"ba"),u'(x"37"),u'(x"b7"),u'(x"00"),u'(x"87"),
u'(x"57"),u'(x"e0"),u'(x"04"),u'(x"77"),u'(x"a9"),u'(x"00"),u'(x"87"),u'(x"57"),u'(x"f0"),u'(x"04"),u'(x"77"),u'(x"9a"),u'(x"00"),u'(x"87"),u'(x"f7"),u'(x"93"),
u'(x"12"),u'(x"f7"),u'(x"8c"),u'(x"74"),u'(x"f7"),u'(x"5c"),u'(x"37"),u'(x"83"),u'(x"c0"),u'(x"6e"),u'(x"37"),u'(x"7b"),u'(x"c1"),u'(x"80"),u'(x"41"),u'(x"a0"),
u'(x"c1"),u'(x"01"),u'(x"62"),u'(x"57"),u'(x"f0"),u'(x"04"),u'(x"f7"),u'(x"01"),u'(x"60"),u'(x"5e"),u'(x"57"),u'(x"e0"),u'(x"04"),u'(x"f7"),u'(x"01"),u'(x"53"),
u'(x"57"),u'(x"f7"),u'(x"22"),u'(x"c0"),u'(x"01"),u'(x"52"),u'(x"c1"),u'(x"80"),u'(x"4f"),u'(x"c1"),u'(x"80"),u'(x"f7"),u'(x"3a"),u'(x"04"),u'(x"f7"),u'(x"35"),
u'(x"01"),u'(x"30"),u'(x"f7"),u'(x"2e"),u'(x"06"),u'(x"f7"),u'(x"29"),u'(x"03"),u'(x"41"),u'(x"a0"),u'(x"02"),u'(x"41"),u'(x"20"),u'(x"c1"),u'(x"39"),u'(x"57"),
u'(x"61"),u'(x"14"),u'(x"57"),u'(x"7a"),u'(x"33"),u'(x"c1"),u'(x"60"),u'(x"57"),u'(x"13"),u'(x"03"),u'(x"b7"),u'(x"8b"),u'(x"08"),u'(x"57"),u'(x"11"),u'(x"05"),
u'(x"37"),u'(x"7f"),u'(x"37"),u'(x"7a"),u'(x"00"),u'(x"1f"),u'(x"57"),u'(x"40"),u'(x"06"),u'(x"57"),u'(x"5b"),u'(x"1c"),u'(x"57"),u'(x"5f"),u'(x"19"),u'(x"c1"),
u'(x"40"),u'(x"13"),u'(x"f7"),u'(x"ce"),u'(x"09"),u'(x"f7"),u'(x"c9"),u'(x"06"),u'(x"f7"),u'(x"c4"),u'(x"03"),u'(x"41"),u'(x"a0"),u'(x"02"),u'(x"41"),u'(x"20"),
u'(x"c1"),u'(x"00"),u'(x"c1"),u'(x"04"),u'(x"00"),u'(x"c0"),u'(x"01"),u'(x"87"),u'(x"00"),u'(x"87"),u'(x"df"),u'(x"70"),u'(x"24"),u'(x"26"),u'(x"66"),u'(x"c1"),
u'(x"72"),u'(x"c0"),u'(x"1e"),u'(x"80"),u'(x"17"),u'(x"80"),u'(x"01"),u'(x"00"),u'(x"37"),u'(x"12"),u'(x"07"),u'(x"b7"),u'(x"06"),u'(x"37"),u'(x"06"),u'(x"c0"),
u'(x"40"),u'(x"48"),u'(x"d7"),u'(x"f8"),u'(x"50"),u'(x"09"),u'(x"f7"),u'(x"f2"),u'(x"06"),u'(x"b7"),u'(x"ec"),u'(x"c0"),u'(x"13"),u'(x"f7"),u'(x"0c"),u'(x"81"),
u'(x"80"),u'(x"df"),u'(x"40"),u'(x"70"),u'(x"02"),u'(x"df"),u'(x"74"),u'(x"fd"),u'(x"1f"),u'(x"76"),u'(x"87"),u'(x"02"),u'(x"df"),u'(x"00"),u'(x"16"),u'(x"26"),
u'(x"66"),u'(x"c0"),u'(x"c2"),u'(x"c1"),u'(x"c0"),u'(x"80"),u'(x"17"),u'(x"20"),u'(x"01"),u'(x"00"),u'(x"01"),u'(x"07"),u'(x"37"),u'(x"ac"),u'(x"c1"),u'(x"02"),
u'(x"c0"),u'(x"c0"),u'(x"48"),u'(x"81"),u'(x"80"),u'(x"df"),u'(x"40"),u'(x"00"),u'(x"02"),u'(x"48"),u'(x"6c"),u'(x"6f"),u'(x"20"),u'(x"6f"),u'(x"6c"),u'(x"3a"),
u'(x"5b"),u'(x"44"),u'(x"32"),u'(x"31"),u'(x"20"),u'(x"74"),u'(x"30"),u'(x"5d"),u'(x"48"),u'(x"6c"),u'(x"6f"),u'(x"20"),u'(x"6f"),u'(x"6c"),u'(x"3a"),u'(x"5b"),
u'(x"44"),u'(x"32"),u'(x"31"),u'(x"20"),u'(x"74"),u'(x"30"),u'(x"5d"),u'(x"3e"),u'(x"5e"),u'(x"f2"),u'(x"fa"),u'(x"02"),u'(x"3a"),u'(x"e2"),u'(x"10"),u'(x"18"),
u'(x"20"),u'(x"28"),u'(x"30"),u'(x"38"),u'(x"40"),u'(x"48"),u'(x"48"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"12"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"10"),u'(x"00"),u'(x"00"),u'(x"10"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),
u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"00"),u'(x"08"),u'(x"18"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"1e"),u'(x"3e"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"62"),u'(x"68"),u'(x"70"),u'(x"00"),u'(x"00"),u'(x"76"),u'(x"80"),u'(x"8a"),u'(x"94"),u'(x"bc"),u'(x"da"),u'(x"dc"),u'(x"de"),
u'(x"00"),u'(x"18"),u'(x"2a"),u'(x"00"),u'(x"42"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"0a"),u'(x"6e"),u'(x"08"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"94"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"30"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"32"),u'(x"00"),u'(x"00"),u'(x"7c"),
u'(x"8c"),u'(x"cc"),u'(x"cc"),u'(x"cc"),u'(x"12"),u'(x"22"),u'(x"2a"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"32"),
u'(x"00"),u'(x"32"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"98"),u'(x"d0"),u'(x"e0"),u'(x"f0"),u'(x"00"),u'(x"28"),u'(x"28"),u'(x"28"),u'(x"10"),
u'(x"28"),u'(x"26"),u'(x"80"),u'(x"e0"),u'(x"34"),u'(x"28"),u'(x"28"),u'(x"8e"),u'(x"28"),u'(x"28"),u'(x"28"),u'(x"28"),u'(x"28"),u'(x"28"),u'(x"28"),u'(x"c2"),
u'(x"28"),u'(x"28"),u'(x"28"),u'(x"28"),u'(x"28"),u'(x"28"),u'(x"28"),u'(x"28"),u'(x"28"),u'(x"28"),u'(x"ee"),u'(x"28"),u'(x"28"),u'(x"08"),u'(x"0e"),u'(x"3c"),
u'(x"28"),u'(x"28"),u'(x"28"),u'(x"ba"),u'(x"46"),u'(x"d6"),u'(x"28"),u'(x"28"),u'(x"28"),u'(x"78"),u'(x"28"),u'(x"28"),u'(x"28"),u'(x"28"),u'(x"28"),u'(x"c6"),
u'(x"24"),u'(x"28"),u'(x"28"),u'(x"28"),u'(x"28"),u'(x"28"),u'(x"28"),u'(x"00"),u'(x"a0"),u'(x"40"),u'(x"e0"),u'(x"80"),u'(x"20"),u'(x"c0"),u'(x"60"),u'(x"00"),
u'(x"a0"),u'(x"40"),u'(x"e0"),u'(x"80"),u'(x"20"),u'(x"c0"),u'(x"60"),u'(x"00"),u'(x"a0"),u'(x"40"),u'(x"e0"),u'(x"80"),u'(x"20"),u'(x"c0"),u'(x"60"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"ff"),u'(x"fe"),u'(x"00"),u'(x"00"),u'(x"e0"),u'(x"60"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"31"),u'(x"00"),u'(x"7a"),u'(x"61"),u'(x"32"),
u'(x"00"),u'(x"78"),u'(x"65"),u'(x"33"),u'(x"00"),u'(x"76"),u'(x"74"),u'(x"35"),u'(x"00"),u'(x"62"),u'(x"67"),u'(x"36"),u'(x"00"),u'(x"6d"),u'(x"75"),u'(x"38"),
u'(x"00"),u'(x"6b"),u'(x"6f"),u'(x"39"),u'(x"00"),u'(x"2f"),u'(x"3b"),u'(x"2d"),u'(x"00"),u'(x"27"),u'(x"5b"),u'(x"00"),u'(x"00"),u'(x"e7"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"7f"),u'(x"00"),u'(x"00"),u'(x"f6"),u'(x"00"),u'(x"ef"),u'(x"f1"),u'(x"f5"),u'(x"1b"),u'(x"00"),u'(x"f2"),u'(x"eb"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"7e"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"21"),u'(x"00"),u'(x"5a"),u'(x"41"),u'(x"40"),
u'(x"00"),u'(x"58"),u'(x"45"),u'(x"23"),u'(x"00"),u'(x"56"),u'(x"54"),u'(x"25"),u'(x"00"),u'(x"42"),u'(x"47"),u'(x"5e"),u'(x"00"),u'(x"4d"),u'(x"55"),u'(x"2a"),
u'(x"00"),u'(x"4b"),u'(x"4f"),u'(x"28"),u'(x"00"),u'(x"3f"),u'(x"3a"),u'(x"5f"),u'(x"00"),u'(x"22"),u'(x"7b"),u'(x"00"),u'(x"00"),u'(x"0d"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"08"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"1b"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"e8"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"ea"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"fa"),u'(x"00"),u'(x"f9"),u'(x"e2"),u'(x"e3"),u'(x"00"),u'(x"00"),u'(x"e5"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00") 
);

signal memo : mem_type := mem_type'(
u'(x"00"),u'(x"01"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"15"),u'(x"02"),u'(x"0a"),u'(x"fe"),u'(x"0a"),u'(x"fe"),u'(x"0a"),u'(x"fe"),u'(x"8a"),u'(x"fe"),u'(x"8a"),u'(x"fe"),u'(x"0a"),
u'(x"fe"),u'(x"0a"),u'(x"fe"),u'(x"15"),u'(x"19"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"1a"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),
u'(x"1a"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"15"),u'(x"00"),u'(x"d0"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"0a"),u'(x"ff"),
u'(x"09"),u'(x"08"),u'(x"15"),u'(x"80"),u'(x"15"),u'(x"00"),u'(x"20"),u'(x"8f"),u'(x"02"),u'(x"15"),u'(x"1a"),u'(x"15"),u'(x"80"),u'(x"25"),u'(x"00"),u'(x"c0"),
u'(x"02"),u'(x"15"),u'(x"1a"),u'(x"94"),u'(x"10"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"8a"),u'(x"fe"),u'(x"8a"),u'(x"fe"),u'(x"8a"),u'(x"fe"),u'(x"8a"),u'(x"fe"),
u'(x"8a"),u'(x"fe"),u'(x"8a"),u'(x"fe"),u'(x"8a"),u'(x"fe"),u'(x"09"),u'(x"14"),u'(x"15"),u'(x"00"),u'(x"fe"),u'(x"15"),u'(x"00"),u'(x"fe"),u'(x"15"),u'(x"00"),
u'(x"fe"),u'(x"15"),u'(x"00"),u'(x"fe"),u'(x"95"),u'(x"00"),u'(x"fe"),u'(x"95"),u'(x"00"),u'(x"fe"),u'(x"95"),u'(x"00"),u'(x"fe"),u'(x"95"),u'(x"00"),u'(x"fe"),
u'(x"15"),u'(x"00"),u'(x"fe"),u'(x"15"),u'(x"00"),u'(x"fe"),u'(x"15"),u'(x"00"),u'(x"fe"),u'(x"8a"),u'(x"fe"),u'(x"8a"),u'(x"fd"),u'(x"8a"),u'(x"fe"),u'(x"95"),
u'(x"00"),u'(x"fe"),u'(x"8a"),u'(x"fe"),u'(x"8a"),u'(x"fe"),u'(x"8a"),u'(x"fe"),u'(x"8a"),u'(x"fe"),u'(x"8a"),u'(x"fd"),u'(x"8a"),u'(x"fd"),u'(x"8a"),u'(x"fe"),
u'(x"8a"),u'(x"fe"),u'(x"8a"),u'(x"fe"),u'(x"8a"),u'(x"fe"),u'(x"8a"),u'(x"fe"),u'(x"0a"),u'(x"c0"),u'(x"0a"),u'(x"c0"),u'(x"0a"),u'(x"c0"),u'(x"0a"),u'(x"c0"),
u'(x"09"),u'(x"0e"),u'(x"10"),u'(x"c0"),u'(x"09"),u'(x"14"),u'(x"0b"),u'(x"03"),u'(x"8a"),u'(x"c0"),u'(x"09"),u'(x"15"),u'(x"0b"),u'(x"03"),u'(x"a0"),u'(x"00"),
u'(x"87"),u'(x"09"),u'(x"03"),u'(x"01"),u'(x"10"),u'(x"09"),u'(x"16"),u'(x"01"),u'(x"09"),u'(x"13"),u'(x"0b"),u'(x"03"),u'(x"8a"),u'(x"c0"),u'(x"45"),u'(x"ff"),
u'(x"09"),u'(x"10"),u'(x"0b"),u'(x"03"),u'(x"9c"),u'(x"1a"),u'(x"0b"),u'(x"03"),u'(x"10"),u'(x"fd"),u'(x"1d"),u'(x"fd"),u'(x"45"),u'(x"ff"),u'(x"65"),u'(x"1a"),
u'(x"12"),u'(x"09"),u'(x"01"),u'(x"a0"),u'(x"00"),u'(x"87"),u'(x"a0"),u'(x"00"),u'(x"82"),u'(x"e5"),u'(x"00"),u'(x"0c"),u'(x"1c"),u'(x"04"),u'(x"10"),u'(x"fd"),
u'(x"0a"),u'(x"fd"),u'(x"01"),u'(x"a0"),u'(x"00"),u'(x"87"),u'(x"a0"),u'(x"00"),u'(x"82"),u'(x"0b"),u'(x"fd"),u'(x"02"),u'(x"10"),u'(x"fd"),u'(x"1d"),u'(x"fd"),
u'(x"20"),u'(x"04"),u'(x"03"),u'(x"20"),u'(x"05"),u'(x"03"),u'(x"01"),u'(x"09"),u'(x"01"),u'(x"45"),u'(x"ff"),u'(x"0c"),u'(x"0c"),u'(x"0c"),u'(x"0c"),u'(x"0c"),
u'(x"45"),u'(x"ff"),u'(x"fd"),u'(x"6d"),u'(x"fd"),u'(x"0a"),u'(x"fd"),u'(x"0b"),u'(x"fd"),u'(x"03"),u'(x"1d"),u'(x"fd"),u'(x"09"),u'(x"01"),u'(x"0a"),u'(x"fd"),
u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"04"),u'(x"04"),u'(x"05"),u'(x"05"),u'(x"05"),u'(x"05"),u'(x"05"),u'(x"05"),u'(x"05"),u'(x"05"),u'(x"06"),u'(x"06"),u'(x"06"),
u'(x"45"),u'(x"ff"),u'(x"8b"),u'(x"fd"),u'(x"02"),u'(x"10"),u'(x"c0"),u'(x"01"),u'(x"10"),u'(x"c0"),u'(x"01"),u'(x"00"),u'(x"35"),u'(x"00"),u'(x"03"),u'(x"55"),
u'(x"00"),u'(x"c0"),u'(x"01"),u'(x"45"),u'(x"00"),u'(x"c0"),u'(x"35"),u'(x"00"),u'(x"03"),u'(x"55"),u'(x"00"),u'(x"c0"),u'(x"01"),u'(x"45"),u'(x"00"),u'(x"c0"),
u'(x"35"),u'(x"00"),u'(x"03"),u'(x"55"),u'(x"00"),u'(x"c0"),u'(x"01"),u'(x"45"),u'(x"00"),u'(x"c0"),u'(x"35"),u'(x"00"),u'(x"03"),u'(x"55"),u'(x"00"),u'(x"c0"),
u'(x"01"),u'(x"45"),u'(x"00"),u'(x"c0"),u'(x"35"),u'(x"00"),u'(x"03"),u'(x"55"),u'(x"00"),u'(x"c0"),u'(x"01"),u'(x"45"),u'(x"00"),u'(x"c0"),u'(x"35"),u'(x"00"),
u'(x"03"),u'(x"55"),u'(x"04"),u'(x"c0"),u'(x"01"),u'(x"45"),u'(x"04"),u'(x"c0"),u'(x"0b"),u'(x"fc"),u'(x"02"),u'(x"35"),u'(x"00"),u'(x"03"),u'(x"55"),u'(x"08"),
u'(x"c0"),u'(x"01"),u'(x"45"),u'(x"08"),u'(x"c0"),u'(x"35"),u'(x"00"),u'(x"03"),u'(x"95"),u'(x"00"),u'(x"fc"),u'(x"01"),u'(x"8a"),u'(x"fc"),u'(x"35"),u'(x"01"),
u'(x"03"),u'(x"55"),u'(x"10"),u'(x"c0"),u'(x"01"),u'(x"45"),u'(x"10"),u'(x"c0"),u'(x"35"),u'(x"02"),u'(x"03"),u'(x"55"),u'(x"20"),u'(x"c0"),u'(x"01"),u'(x"45"),
u'(x"20"),u'(x"c0"),u'(x"00"),u'(x"1d"),u'(x"fc"),u'(x"0c"),u'(x"45"),u'(x"fc"),u'(x"55"),u'(x"90"),u'(x"90"),u'(x"35"),u'(x"20"),u'(x"c0"),u'(x"02"),u'(x"0a"),
u'(x"fc"),u'(x"45"),u'(x"fe"),u'(x"fc"),u'(x"1d"),u'(x"fc"),u'(x"c0"),u'(x"00"),u'(x"25"),u'(x"01"),u'(x"87"),u'(x"0c"),u'(x"45"),u'(x"fc"),u'(x"55"),u'(x"90"),
u'(x"c5"),u'(x"00"),u'(x"01"),u'(x"45"),u'(x"fe"),u'(x"0c"),u'(x"45"),u'(x"fc"),u'(x"55"),u'(x"90"),u'(x"d5"),u'(x"00"),u'(x"01"),u'(x"00"),u'(x"25"),u'(x"01"),
u'(x"87"),u'(x"0c"),u'(x"45"),u'(x"fc"),u'(x"55"),u'(x"90"),u'(x"c5"),u'(x"00"),u'(x"01"),u'(x"45"),u'(x"fe"),u'(x"0c"),u'(x"45"),u'(x"fc"),u'(x"55"),u'(x"90"),
u'(x"d5"),u'(x"00"),u'(x"01"),u'(x"00"),u'(x"00"),u'(x"10"),u'(x"fb"),u'(x"10"),u'(x"c0"),u'(x"00"),u'(x"35"),u'(x"00"),u'(x"03"),u'(x"55"),u'(x"00"),u'(x"c0"),
u'(x"01"),u'(x"45"),u'(x"00"),u'(x"c0"),u'(x"35"),u'(x"00"),u'(x"03"),u'(x"55"),u'(x"00"),u'(x"c0"),u'(x"01"),u'(x"45"),u'(x"00"),u'(x"c0"),u'(x"35"),u'(x"00"),
u'(x"03"),u'(x"55"),u'(x"01"),u'(x"c0"),u'(x"01"),u'(x"45"),u'(x"01"),u'(x"c0"),u'(x"35"),u'(x"00"),u'(x"03"),u'(x"55"),u'(x"02"),u'(x"c0"),u'(x"01"),u'(x"45"),
u'(x"02"),u'(x"c0"),u'(x"35"),u'(x"00"),u'(x"03"),u'(x"09"),u'(x"11"),u'(x"0b"),u'(x"fb"),u'(x"02"),u'(x"35"),u'(x"00"),u'(x"03"),u'(x"55"),u'(x"80"),u'(x"c0"),
u'(x"01"),u'(x"45"),u'(x"80"),u'(x"c0"),u'(x"00"),u'(x"1d"),u'(x"fb"),u'(x"0c"),u'(x"45"),u'(x"fc"),u'(x"55"),u'(x"94"),u'(x"90"),u'(x"0a"),u'(x"fb"),u'(x"45"),
u'(x"fe"),u'(x"fb"),u'(x"1d"),u'(x"fb"),u'(x"c0"),u'(x"00"),u'(x"25"),u'(x"01"),u'(x"87"),u'(x"0c"),u'(x"45"),u'(x"fc"),u'(x"55"),u'(x"90"),u'(x"c5"),u'(x"00"),
u'(x"01"),u'(x"45"),u'(x"fe"),u'(x"0c"),u'(x"45"),u'(x"fc"),u'(x"55"),u'(x"90"),u'(x"d5"),u'(x"00"),u'(x"01"),u'(x"00"),u'(x"25"),u'(x"01"),u'(x"87"),u'(x"0c"),
u'(x"45"),u'(x"fc"),u'(x"55"),u'(x"90"),u'(x"c5"),u'(x"00"),u'(x"01"),u'(x"45"),u'(x"fe"),u'(x"0c"),u'(x"45"),u'(x"fc"),u'(x"55"),u'(x"90"),u'(x"d5"),u'(x"00"),
u'(x"01"),u'(x"00"),u'(x"45"),u'(x"ff"),u'(x"e5"),u'(x"00"),u'(x"45"),u'(x"ff"),u'(x"0c"),u'(x"1c"),u'(x"09"),u'(x"09"),u'(x"00"),u'(x"09"),u'(x"02"),u'(x"15"),
u'(x"00"),u'(x"09"),u'(x"13"),u'(x"00"),u'(x"09"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"13"),u'(x"00"),u'(x"09"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"09"),
u'(x"13"),u'(x"00"),u'(x"09"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"13"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"09"),
u'(x"13"),u'(x"0a"),u'(x"02"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"12"),u'(x"0a"),u'(x"02"),u'(x"00"),u'(x"15"),
u'(x"00"),u'(x"09"),u'(x"12"),u'(x"0b"),u'(x"fa"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"12"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"12"),u'(x"8b"),
u'(x"fa"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"12"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"12"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"12"),u'(x"8b"),
u'(x"f9"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"12"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"12"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"12"),u'(x"8b"),
u'(x"f9"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"12"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"12"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"12"),u'(x"8b"),
u'(x"f9"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"12"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"12"),u'(x"00"),u'(x"8b"),u'(x"f9"),u'(x"02"),u'(x"15"),u'(x"00"),
u'(x"09"),u'(x"12"),u'(x"00"),u'(x"00"),u'(x"8b"),u'(x"f9"),u'(x"02"),u'(x"09"),u'(x"ff"),u'(x"00"),u'(x"09"),u'(x"01"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"12"),
u'(x"00"),u'(x"8b"),u'(x"f9"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"12"),u'(x"00"),u'(x"09"),u'(x"01"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"12"),u'(x"00"),
u'(x"8b"),u'(x"f9"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"11"),u'(x"00"),u'(x"09"),u'(x"01"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"11"),u'(x"00"),u'(x"8b"),
u'(x"f9"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"11"),u'(x"00"),u'(x"09"),u'(x"01"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"11"),u'(x"00"),u'(x"8b"),u'(x"f9"),
u'(x"02"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"11"),u'(x"00"),u'(x"09"),u'(x"01"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"11"),u'(x"00"),u'(x"8b"),u'(x"f9"),u'(x"02"),
u'(x"15"),u'(x"00"),u'(x"09"),u'(x"11"),u'(x"00"),u'(x"09"),u'(x"01"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"11"),u'(x"00"),u'(x"8b"),u'(x"f8"),u'(x"02"),u'(x"15"),
u'(x"00"),u'(x"09"),u'(x"11"),u'(x"00"),u'(x"09"),u'(x"01"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"11"),u'(x"00"),u'(x"8b"),u'(x"f8"),u'(x"02"),u'(x"15"),u'(x"00"),
u'(x"09"),u'(x"11"),u'(x"00"),u'(x"09"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"11"),u'(x"00"),u'(x"8b"),u'(x"f8"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"09"),
u'(x"11"),u'(x"00"),u'(x"09"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"11"),u'(x"00"),u'(x"8b"),u'(x"f8"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"11"),
u'(x"00"),u'(x"09"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"11"),u'(x"00"),u'(x"8b"),u'(x"f8"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"11"),u'(x"00"),
u'(x"09"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"10"),u'(x"00"),u'(x"8b"),u'(x"f8"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"10"),u'(x"00"),u'(x"09"),
u'(x"00"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"10"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"10"),u'(x"00"),u'(x"00"),u'(x"09"),u'(x"00"),
u'(x"15"),u'(x"00"),u'(x"09"),u'(x"10"),u'(x"00"),u'(x"09"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"10"),u'(x"00"),u'(x"09"),u'(x"00"),u'(x"15"),u'(x"00"),
u'(x"09"),u'(x"10"),u'(x"00"),u'(x"09"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"10"),u'(x"00"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"10"),u'(x"8b"),
u'(x"f7"),u'(x"02"),u'(x"8b"),u'(x"f7"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"10"),u'(x"01"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"10"),u'(x"01"),u'(x"00"),
u'(x"15"),u'(x"00"),u'(x"09"),u'(x"10"),u'(x"8b"),u'(x"f7"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"10"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"10"),
u'(x"00"),u'(x"09"),u'(x"06"),u'(x"06"),u'(x"06"),u'(x"06"),u'(x"06"),u'(x"07"),u'(x"07"),u'(x"07"),u'(x"07"),u'(x"07"),u'(x"07"),u'(x"07"),u'(x"07"),u'(x"07"),
u'(x"08"),u'(x"08"),u'(x"08"),u'(x"08"),u'(x"08"),u'(x"08"),u'(x"08"),u'(x"08"),u'(x"08"),u'(x"09"),u'(x"09"),u'(x"09"),u'(x"09"),u'(x"09"),u'(x"09"),u'(x"09"),
u'(x"09"),u'(x"09"),u'(x"00"),u'(x"15"),u'(x"80"),u'(x"15"),u'(x"8f"),u'(x"15"),u'(x"00"),u'(x"20"),u'(x"87"),u'(x"00"),u'(x"1d"),u'(x"f6"),u'(x"0a"),u'(x"95"),
u'(x"00"),u'(x"c0"),u'(x"09"),u'(x"00"),u'(x"00"),u'(x"1d"),u'(x"f6"),u'(x"0a"),u'(x"95"),u'(x"00"),u'(x"c0"),u'(x"09"),u'(x"00"),u'(x"00"),u'(x"1d"),u'(x"f6"),
u'(x"0a"),u'(x"95"),u'(x"00"),u'(x"c0"),u'(x"09"),u'(x"00"),u'(x"00"),u'(x"1d"),u'(x"f6"),u'(x"0a"),u'(x"8a"),u'(x"c0"),u'(x"00"),u'(x"2d"),u'(x"f6"),u'(x"00"),
u'(x"83"),u'(x"15"),u'(x"00"),u'(x"f6"),u'(x"1d"),u'(x"f6"),u'(x"10"),u'(x"0a"),u'(x"0c"),u'(x"1c"),u'(x"1d"),u'(x"65"),u'(x"00"),u'(x"0c"),u'(x"1c"),u'(x"1d"),
u'(x"15"),u'(x"00"),u'(x"20"),u'(x"87"),u'(x"00"),u'(x"10"),u'(x"10"),u'(x"15"),u'(x"c0"),u'(x"15"),u'(x"c0"),u'(x"0a"),u'(x"20"),u'(x"87"),u'(x"15"),u'(x"15"),
u'(x"00"),u'(x"10"),u'(x"10"),u'(x"15"),u'(x"c0"),u'(x"6d"),u'(x"f6"),u'(x"0a"),u'(x"15"),u'(x"c0"),u'(x"8a"),u'(x"20"),u'(x"87"),u'(x"15"),u'(x"15"),u'(x"00"),
u'(x"10"),u'(x"10"),u'(x"15"),u'(x"c0"),u'(x"10"),u'(x"6d"),u'(x"f6"),u'(x"8a"),u'(x"20"),u'(x"87"),u'(x"15"),u'(x"15"),u'(x"00"),u'(x"10"),u'(x"10"),u'(x"15"),
u'(x"80"),u'(x"15"),u'(x"8f"),u'(x"15"),u'(x"00"),u'(x"20"),u'(x"87"),u'(x"15"),u'(x"00"),u'(x"f5"),u'(x"15"),u'(x"00"),u'(x"f5"),u'(x"8a"),u'(x"f5"),u'(x"09"),
u'(x"ff"),u'(x"15"),u'(x"15"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"c0"),u'(x"02"),u'(x"95"),u'(x"00"),u'(x"f6"),u'(x"00"),u'(x"8a"),u'(x"f6"),u'(x"00"),u'(x"1d"),
u'(x"f5"),u'(x"f5"),u'(x"1d"),u'(x"f5"),u'(x"f5"),u'(x"9d"),u'(x"f5"),u'(x"f5"),u'(x"9d"),u'(x"f5"),u'(x"f5"),u'(x"9d"),u'(x"f5"),u'(x"f5"),u'(x"00"),u'(x"1d"),
u'(x"f5"),u'(x"f5"),u'(x"1d"),u'(x"f5"),u'(x"f5"),u'(x"9d"),u'(x"f5"),u'(x"f5"),u'(x"9d"),u'(x"f5"),u'(x"f5"),u'(x"9d"),u'(x"f5"),u'(x"f5"),u'(x"09"),u'(x"06"),
u'(x"00"),u'(x"8a"),u'(x"f5"),u'(x"00"),u'(x"95"),u'(x"00"),u'(x"f5"),u'(x"00"),u'(x"8a"),u'(x"f5"),u'(x"00"),u'(x"0a"),u'(x"f5"),u'(x"09"),u'(x"06"),u'(x"00"),
u'(x"0a"),u'(x"f5"),u'(x"09"),u'(x"06"),u'(x"00"),u'(x"0a"),u'(x"f5"),u'(x"09"),u'(x"06"),u'(x"00"),u'(x"8b"),u'(x"f5"),u'(x"02"),u'(x"2d"),u'(x"f5"),u'(x"f5"),
u'(x"03"),u'(x"0a"),u'(x"f5"),u'(x"01"),u'(x"09"),u'(x"06"),u'(x"8a"),u'(x"f5"),u'(x"00"),u'(x"0a"),u'(x"f5"),u'(x"09"),u'(x"06"),u'(x"00"),u'(x"15"),u'(x"00"),
u'(x"f5"),u'(x"2d"),u'(x"f5"),u'(x"f5"),u'(x"03"),u'(x"0a"),u'(x"f5"),u'(x"01"),u'(x"09"),u'(x"06"),u'(x"8a"),u'(x"f5"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"8b"),
u'(x"f5"),u'(x"02"),u'(x"1d"),u'(x"f5"),u'(x"0a"),u'(x"95"),u'(x"00"),u'(x"01"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"f4"),u'(x"15"),u'(x"00"),u'(x"f4"),u'(x"00"),
u'(x"25"),u'(x"00"),u'(x"f4"),u'(x"03"),u'(x"0a"),u'(x"f4"),u'(x"01"),u'(x"09"),u'(x"06"),u'(x"8a"),u'(x"f4"),u'(x"00"),u'(x"09"),u'(x"06"),u'(x"15"),u'(x"8f"),
u'(x"15"),u'(x"00"),u'(x"20"),u'(x"87"),u'(x"00"),u'(x"09"),u'(x"05"),u'(x"1d"),u'(x"f4"),u'(x"0c"),u'(x"1c"),u'(x"1d"),u'(x"15"),u'(x"00"),u'(x"20"),u'(x"87"),
u'(x"00"),u'(x"8b"),u'(x"f5"),u'(x"02"),u'(x"2d"),u'(x"f4"),u'(x"f4"),u'(x"03"),u'(x"0a"),u'(x"f4"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"f4"),u'(x"03"),u'(x"0a"),
u'(x"f4"),u'(x"01"),u'(x"09"),u'(x"06"),u'(x"8a"),u'(x"f4"),u'(x"00"),u'(x"8b"),u'(x"f4"),u'(x"02"),u'(x"09"),u'(x"02"),u'(x"00"),u'(x"95"),u'(x"00"),u'(x"09"),
u'(x"0d"),u'(x"95"),u'(x"00"),u'(x"09"),u'(x"0d"),u'(x"95"),u'(x"00"),u'(x"09"),u'(x"0d"),u'(x"00"),u'(x"00"),u'(x"f5"),u'(x"10"),u'(x"09"),u'(x"05"),u'(x"10"),
u'(x"1d"),u'(x"f4"),u'(x"0c"),u'(x"1c"),u'(x"1d"),u'(x"10"),u'(x"0a"),u'(x"0a"),u'(x"20"),u'(x"03"),u'(x"18"),u'(x"20"),u'(x"82"),u'(x"15"),u'(x"00"),u'(x"25"),
u'(x"00"),u'(x"f4"),u'(x"03"),u'(x"0a"),u'(x"f4"),u'(x"01"),u'(x"15"),u'(x"00"),u'(x"ed"),u'(x"f4"),u'(x"f4"),u'(x"09"),u'(x"05"),u'(x"8a"),u'(x"f4"),u'(x"00"),
u'(x"6d"),u'(x"f4"),u'(x"f4"),u'(x"09"),u'(x"05"),u'(x"8a"),u'(x"f4"),u'(x"00"),u'(x"6d"),u'(x"f4"),u'(x"f3"),u'(x"09"),u'(x"05"),u'(x"8a"),u'(x"f3"),u'(x"00"),
u'(x"ed"),u'(x"f4"),u'(x"f3"),u'(x"09"),u'(x"05"),u'(x"8a"),u'(x"f3"),u'(x"00"),u'(x"1d"),u'(x"f4"),u'(x"f3"),u'(x"1d"),u'(x"f4"),u'(x"f3"),u'(x"09"),u'(x"05"),
u'(x"8a"),u'(x"f3"),u'(x"00"),u'(x"09"),u'(x"05"),u'(x"0b"),u'(x"f4"),u'(x"02"),u'(x"09"),u'(x"fd"),u'(x"15"),u'(x"8f"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"f4"),
u'(x"02"),u'(x"09"),u'(x"fd"),u'(x"10"),u'(x"0a"),u'(x"15"),u'(x"80"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"f4"),u'(x"03"),u'(x"25"),u'(x"00"),u'(x"f4"),u'(x"03"),
u'(x"01"),u'(x"09"),u'(x"fd"),u'(x"15"),u'(x"80"),u'(x"15"),u'(x"8f"),u'(x"01"),u'(x"15"),u'(x"00"),u'(x"20"),u'(x"87"),u'(x"01"),u'(x"8a"),u'(x"f3"),u'(x"00"),
u'(x"09"),u'(x"04"),u'(x"0b"),u'(x"f3"),u'(x"02"),u'(x"1d"),u'(x"f3"),u'(x"0c"),u'(x"1c"),u'(x"1d"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"f3"),u'(x"02"),u'(x"10"),
u'(x"0a"),u'(x"1d"),u'(x"f3"),u'(x"0a"),u'(x"0c"),u'(x"1c"),u'(x"1d"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"f3"),u'(x"02"),u'(x"1d"),u'(x"f3"),u'(x"0a"),u'(x"0c"),
u'(x"1c"),u'(x"1d"),u'(x"1d"),u'(x"f3"),u'(x"0c"),u'(x"1c"),u'(x"1d"),u'(x"01"),u'(x"15"),u'(x"00"),u'(x"20"),u'(x"87"),u'(x"01"),u'(x"8a"),u'(x"f3"),u'(x"00"),
u'(x"10"),u'(x"2d"),u'(x"f3"),u'(x"f3"),u'(x"82"),u'(x"1d"),u'(x"f3"),u'(x"0c"),u'(x"1c"),u'(x"1d"),u'(x"1d"),u'(x"f3"),u'(x"ed"),u'(x"f3"),u'(x"0c"),u'(x"1c"),
u'(x"1d"),u'(x"1d"),u'(x"f2"),u'(x"0a"),u'(x"6d"),u'(x"f2"),u'(x"0a"),u'(x"0c"),u'(x"1c"),u'(x"1d"),u'(x"20"),u'(x"83"),u'(x"18"),u'(x"20"),u'(x"82"),u'(x"0a"),
u'(x"0a"),u'(x"95"),u'(x"00"),u'(x"20"),u'(x"82"),u'(x"15"),u'(x"00"),u'(x"f2"),u'(x"15"),u'(x"00"),u'(x"10"),u'(x"2d"),u'(x"f2"),u'(x"f2"),u'(x"82"),u'(x"1d"),
u'(x"f2"),u'(x"6d"),u'(x"f2"),u'(x"0a"),u'(x"0a"),u'(x"10"),u'(x"6d"),u'(x"f3"),u'(x"1d"),u'(x"f2"),u'(x"ed"),u'(x"f2"),u'(x"20"),u'(x"86"),u'(x"10"),u'(x"0c"),
u'(x"0c"),u'(x"1c"),u'(x"1d"),u'(x"1c"),u'(x"1d"),u'(x"1d"),u'(x"f2"),u'(x"0c"),u'(x"1c"),u'(x"1d"),u'(x"14"),u'(x"20"),u'(x"87"),u'(x"95"),u'(x"00"),u'(x"0a"),
u'(x"20"),u'(x"87"),u'(x"15"),u'(x"00"),u'(x"f2"),u'(x"15"),u'(x"00"),u'(x"10"),u'(x"1d"),u'(x"f2"),u'(x"0c"),u'(x"1c"),u'(x"1d"),u'(x"09"),u'(x"03"),u'(x"10"),
u'(x"6d"),u'(x"f2"),u'(x"6d"),u'(x"f2"),u'(x"20"),u'(x"87"),u'(x"10"),u'(x"01"),u'(x"14"),u'(x"20"),u'(x"87"),u'(x"15"),u'(x"00"),u'(x"20"),u'(x"87"),u'(x"15"),
u'(x"00"),u'(x"10"),u'(x"1d"),u'(x"f2"),u'(x"0c"),u'(x"1c"),u'(x"1d"),u'(x"09"),u'(x"03"),u'(x"10"),u'(x"6d"),u'(x"f2"),u'(x"6d"),u'(x"f2"),u'(x"20"),u'(x"87"),
u'(x"10"),u'(x"15"),u'(x"00"),u'(x"20"),u'(x"87"),u'(x"15"),u'(x"00"),u'(x"15"),u'(x"0f"),u'(x"94"),u'(x"09"),u'(x"0b"),u'(x"20"),u'(x"0f"),u'(x"02"),u'(x"00"),
u'(x"5b"),u'(x"31"),u'(x"36"),u'(x"00"),u'(x"09"),u'(x"fe"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"f2"),u'(x"02"),u'(x"1d"),u'(x"f1"),u'(x"0a"),u'(x"8a"),u'(x"01"),
u'(x"01"),u'(x"25"),u'(x"00"),u'(x"f2"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"0a"),u'(x"8a"),u'(x"01"),u'(x"0a"),u'(x"0b"),u'(x"02"),u'(x"00"),u'(x"0a"),u'(x"20"),
u'(x"f2"),u'(x"82"),u'(x"1c"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"02"),u'(x"95"),u'(x"00"),u'(x"f2"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"02"),u'(x"95"),u'(x"00"),
u'(x"f2"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"02"),u'(x"95"),u'(x"00"),u'(x"f1"),u'(x"09"),u'(x"fb"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"02"),u'(x"95"),u'(x"00"),
u'(x"f1"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"02"),u'(x"95"),u'(x"00"),u'(x"f1"),u'(x"8a"),u'(x"f1"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"02"),u'(x"95"),u'(x"00"),
u'(x"f1"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"02"),u'(x"45"),u'(x"00"),u'(x"c0"),u'(x"01"),u'(x"0a"),u'(x"0a"),u'(x"01"),u'(x"00"),u'(x"0a"),u'(x"20"),u'(x"f1"),
u'(x"82"),u'(x"1c"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"02"),u'(x"95"),u'(x"00"),u'(x"f1"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"02"),u'(x"95"),u'(x"00"),u'(x"f1"),
u'(x"01"),u'(x"25"),u'(x"00"),u'(x"02"),u'(x"95"),u'(x"00"),u'(x"f1"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"02"),u'(x"95"),u'(x"00"),u'(x"f1"),u'(x"09"),u'(x"fa"),
u'(x"01"),u'(x"25"),u'(x"00"),u'(x"02"),u'(x"95"),u'(x"00"),u'(x"f1"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"02"),u'(x"95"),u'(x"00"),u'(x"f1"),u'(x"8a"),u'(x"f0"),
u'(x"01"),u'(x"25"),u'(x"00"),u'(x"02"),u'(x"95"),u'(x"00"),u'(x"f1"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"02"),u'(x"55"),u'(x"00"),u'(x"c0"),u'(x"01"),u'(x"0a"),
u'(x"0a"),u'(x"01"),u'(x"00"),u'(x"0a"),u'(x"20"),u'(x"f1"),u'(x"82"),u'(x"1c"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"02"),u'(x"8a"),u'(x"f0"),u'(x"01"),u'(x"25"),
u'(x"00"),u'(x"02"),u'(x"d5"),u'(x"00"),u'(x"f0"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"02"),u'(x"d5"),u'(x"00"),u'(x"f0"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"02"),
u'(x"d5"),u'(x"00"),u'(x"f0"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"02"),u'(x"d5"),u'(x"00"),u'(x"f0"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"02"),u'(x"c5"),u'(x"00"),
u'(x"f0"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"02"),u'(x"c5"),u'(x"00"),u'(x"f0"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"02"),u'(x"c5"),u'(x"00"),u'(x"f0"),u'(x"01"),
u'(x"25"),u'(x"00"),u'(x"02"),u'(x"c5"),u'(x"00"),u'(x"f0"),u'(x"01"),u'(x"0a"),u'(x"0a"),u'(x"01"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"f0"),u'(x"03"),u'(x"25"),
u'(x"00"),u'(x"f0"),u'(x"03"),u'(x"01"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"09"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"09"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"09"),
u'(x"15"),u'(x"00"),u'(x"09"),u'(x"09"),u'(x"01"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"08"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"08"),u'(x"1d"),u'(x"ef"),u'(x"0a"),
u'(x"0a"),u'(x"0a"),u'(x"e5"),u'(x"00"),u'(x"80"),u'(x"65"),u'(x"00"),u'(x"0b"),u'(x"03"),u'(x"65"),u'(x"00"),u'(x"09"),u'(x"08"),u'(x"10"),u'(x"09"),u'(x"08"),
u'(x"15"),u'(x"00"),u'(x"09"),u'(x"08"),u'(x"1d"),u'(x"ef"),u'(x"0a"),u'(x"0a"),u'(x"0a"),u'(x"e5"),u'(x"00"),u'(x"80"),u'(x"65"),u'(x"00"),u'(x"0b"),u'(x"03"),
u'(x"65"),u'(x"00"),u'(x"09"),u'(x"08"),u'(x"10"),u'(x"09"),u'(x"08"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"08"),u'(x"00"),u'(x"1d"),u'(x"ef"),u'(x"0b"),u'(x"03"),
u'(x"1d"),u'(x"ef"),u'(x"0b"),u'(x"03"),u'(x"20"),u'(x"86"),u'(x"10"),u'(x"ef"),u'(x"10"),u'(x"ef"),u'(x"e0"),u'(x"0a"),u'(x"10"),u'(x"ef"),u'(x"01"),u'(x"15"),
u'(x"00"),u'(x"ef"),u'(x"15"),u'(x"00"),u'(x"ef"),u'(x"15"),u'(x"00"),u'(x"ef"),u'(x"15"),u'(x"00"),u'(x"10"),u'(x"ef"),u'(x"10"),u'(x"ef"),u'(x"09"),u'(x"00"),
u'(x"8a"),u'(x"ef"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"ef"),u'(x"02"),u'(x"15"),u'(x"12"),u'(x"94"),u'(x"09"),u'(x"08"),u'(x"20"),u'(x"12"),u'(x"02"),u'(x"01"),
u'(x"25"),u'(x"00"),u'(x"ef"),u'(x"02"),u'(x"15"),u'(x"11"),u'(x"94"),u'(x"09"),u'(x"08"),u'(x"20"),u'(x"12"),u'(x"02"),u'(x"01"),u'(x"00"),u'(x"5b"),u'(x"3b"),
u'(x"3b"),u'(x"3b"),u'(x"31"),u'(x"3b"),u'(x"31"),u'(x"3b"),u'(x"3b"),u'(x"78"),u'(x"5b"),u'(x"3b"),u'(x"3b"),u'(x"3b"),u'(x"31"),u'(x"3b"),u'(x"31"),u'(x"3b"),
u'(x"3b"),u'(x"78"),u'(x"00"),u'(x"ef"),u'(x"00"),u'(x"10"),u'(x"2d"),u'(x"ee"),u'(x"00"),u'(x"04"),u'(x"15"),u'(x"00"),u'(x"ee"),u'(x"2d"),u'(x"ee"),u'(x"00"),
u'(x"07"),u'(x"15"),u'(x"00"),u'(x"ee"),u'(x"1d"),u'(x"ee"),u'(x"20"),u'(x"00"),u'(x"04"),u'(x"15"),u'(x"00"),u'(x"ee"),u'(x"01"),u'(x"20"),u'(x"00"),u'(x"07"),
u'(x"15"),u'(x"00"),u'(x"ee"),u'(x"01"),u'(x"8b"),u'(x"ee"),u'(x"03"),u'(x"20"),u'(x"ee"),u'(x"07"),u'(x"1d"),u'(x"ee"),u'(x"10"),u'(x"ee"),u'(x"6d"),u'(x"ee"),
u'(x"0a"),u'(x"0a"),u'(x"0c"),u'(x"1c"),u'(x"1d"),u'(x"1d"),u'(x"ee"),u'(x"0a"),u'(x"0c"),u'(x"60"),u'(x"15"),u'(x"00"),u'(x"10"),u'(x"10"),u'(x"10"),u'(x"1d"),
u'(x"ee"),u'(x"10"),u'(x"0a"),u'(x"0c"),u'(x"0c"),u'(x"1c"),u'(x"1d"),u'(x"1c"),u'(x"1d"),u'(x"1d"),u'(x"ee"),u'(x"0c"),u'(x"1c"),u'(x"1d"),u'(x"14"),u'(x"20"),
u'(x"87"),u'(x"15"),u'(x"00"),u'(x"20"),u'(x"87"),u'(x"1d"),u'(x"ee"),u'(x"10"),u'(x"0a"),u'(x"65"),u'(x"c0"),u'(x"65"),u'(x"c0"),u'(x"1d"),u'(x"ee"),u'(x"65"),
u'(x"c0"),u'(x"94"),u'(x"20"),u'(x"87"),u'(x"8a"),u'(x"15"),u'(x"15"),u'(x"15"),u'(x"00"),u'(x"10"),u'(x"10"),u'(x"10"),u'(x"1d"),u'(x"ee"),u'(x"10"),u'(x"0a"),
u'(x"0c"),u'(x"0c"),u'(x"1c"),u'(x"1d"),u'(x"1c"),u'(x"1d"),u'(x"1d"),u'(x"ed"),u'(x"0a"),u'(x"0c"),u'(x"1c"),u'(x"1d"),u'(x"18"),u'(x"20"),u'(x"82"),u'(x"15"),
u'(x"00"),u'(x"20"),u'(x"82"),u'(x"1d"),u'(x"ed"),u'(x"10"),u'(x"0a"),u'(x"65"),u'(x"c0"),u'(x"65"),u'(x"c0"),u'(x"1d"),u'(x"ed"),u'(x"0a"),u'(x"65"),u'(x"c0"),
u'(x"98"),u'(x"20"),u'(x"82"),u'(x"8a"),u'(x"15"),u'(x"15"),u'(x"15"),u'(x"00"),u'(x"8b"),u'(x"ed"),u'(x"03"),u'(x"8b"),u'(x"ed"),u'(x"02"),u'(x"2d"),u'(x"ed"),
u'(x"00"),u'(x"02"),u'(x"2d"),u'(x"ed"),u'(x"ed"),u'(x"86"),u'(x"15"),u'(x"00"),u'(x"ed"),u'(x"65"),u'(x"00"),u'(x"ed"),u'(x"01"),u'(x"09"),u'(x"ff"),u'(x"15"),
u'(x"00"),u'(x"ed"),u'(x"8a"),u'(x"ed"),u'(x"09"),u'(x"fe"),u'(x"00"),u'(x"09"),u'(x"ff"),u'(x"ad"),u'(x"ed"),u'(x"00"),u'(x"02"),u'(x"20"),u'(x"00"),u'(x"87"),
u'(x"20"),u'(x"00"),u'(x"03"),u'(x"e5"),u'(x"00"),u'(x"01"),u'(x"ad"),u'(x"ed"),u'(x"00"),u'(x"02"),u'(x"20"),u'(x"00"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"01"),
u'(x"8b"),u'(x"ed"),u'(x"03"),u'(x"10"),u'(x"10"),u'(x"10"),u'(x"10"),u'(x"1d"),u'(x"ed"),u'(x"0c"),u'(x"1c"),u'(x"1d"),u'(x"10"),u'(x"0a"),u'(x"0a"),u'(x"20"),
u'(x"03"),u'(x"18"),u'(x"20"),u'(x"82"),u'(x"15"),u'(x"15"),u'(x"15"),u'(x"90"),u'(x"9d"),u'(x"ed"),u'(x"0a"),u'(x"2d"),u'(x"ec"),u'(x"00"),u'(x"03"),u'(x"87"),
u'(x"8b"),u'(x"ed"),u'(x"03"),u'(x"95"),u'(x"00"),u'(x"ec"),u'(x"01"),u'(x"65"),u'(x"00"),u'(x"ec"),u'(x"01"),u'(x"00"),u'(x"20"),u'(x"00"),u'(x"86"),u'(x"10"),
u'(x"0c"),u'(x"1c"),u'(x"1c"),u'(x"0b"),u'(x"03"),u'(x"09"),u'(x"0a"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"25"),u'(x"00"),u'(x"c0"),u'(x"03"),u'(x"15"),u'(x"14"),
u'(x"94"),u'(x"09"),u'(x"05"),u'(x"20"),u'(x"14"),u'(x"02"),u'(x"00"),u'(x"15"),u'(x"14"),u'(x"94"),u'(x"09"),u'(x"05"),u'(x"20"),u'(x"14"),u'(x"02"),u'(x"00"),
u'(x"74"),u'(x"30"),u'(x"5b"),u'(x"64"),u'(x"32"),u'(x"31"),u'(x"5d"),u'(x"74"),u'(x"30"),u'(x"5b"),u'(x"64"),u'(x"32"),u'(x"31"),u'(x"5d"),u'(x"e5"),u'(x"00"),
u'(x"ec"),u'(x"09"),u'(x"fd"),u'(x"8a"),u'(x"ec"),u'(x"00"),u'(x"1d"),u'(x"ec"),u'(x"15"),u'(x"01"),u'(x"60"),u'(x"0a"),u'(x"1d"),u'(x"ec"),u'(x"0a"),u'(x"9c"),
u'(x"c0"),u'(x"8b"),u'(x"03"),u'(x"25"),u'(x"00"),u'(x"ec"),u'(x"03"),u'(x"01"),u'(x"25"),u'(x"00"),u'(x"ec"),u'(x"03"),u'(x"0a"),u'(x"ec"),u'(x"0a"),u'(x"8b"),
u'(x"03"),u'(x"09"),u'(x"fd"),u'(x"8a"),u'(x"ec"),u'(x"00"),u'(x"8b"),u'(x"ec"),u'(x"03"),u'(x"15"),u'(x"00"),u'(x"ec"),u'(x"8b"),u'(x"ec"),u'(x"03"),u'(x"2d"),
u'(x"ec"),u'(x"ec"),u'(x"87"),u'(x"09"),u'(x"fd"),u'(x"01"),u'(x"2d"),u'(x"eb"),u'(x"ec"),u'(x"87"),u'(x"2d"),u'(x"eb"),u'(x"ec"),u'(x"82"),u'(x"02"),u'(x"09"),
u'(x"fd"),u'(x"01"),u'(x"65"),u'(x"00"),u'(x"eb"),u'(x"01"),u'(x"8a"),u'(x"eb"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"eb"),u'(x"09"),u'(x"fd"),u'(x"8a"),u'(x"eb"),
u'(x"00"),u'(x"9d"),u'(x"eb"),u'(x"eb"),u'(x"00"),u'(x"9d"),u'(x"eb"),u'(x"eb"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ec"),u'(x"8a"),u'(x"eb"),u'(x"00"),u'(x"8b"),
u'(x"ec"),u'(x"03"),u'(x"09"),u'(x"ee"),u'(x"01"),u'(x"a0"),u'(x"00"),u'(x"87"),u'(x"a0"),u'(x"00"),u'(x"86"),u'(x"09"),u'(x"fe"),u'(x"01"),u'(x"00"),u'(x"a0"),
u'(x"00"),u'(x"87"),u'(x"a0"),u'(x"00"),u'(x"86"),u'(x"45"),u'(x"ff"),u'(x"0c"),u'(x"65"),u'(x"1c"),u'(x"12"),u'(x"1d"),u'(x"eb"),u'(x"ec"),u'(x"0b"),u'(x"ec"),
u'(x"02"),u'(x"15"),u'(x"00"),u'(x"eb"),u'(x"1d"),u'(x"eb"),u'(x"eb"),u'(x"0b"),u'(x"eb"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"eb"),u'(x"09"),u'(x"15"),u'(x"00"),
u'(x"eb"),u'(x"01"),u'(x"a0"),u'(x"00"),u'(x"87"),u'(x"a0"),u'(x"00"),u'(x"82"),u'(x"1d"),u'(x"eb"),u'(x"20"),u'(x"00"),u'(x"87"),u'(x"15"),u'(x"00"),u'(x"1c"),
u'(x"01"),u'(x"0c"),u'(x"0c"),u'(x"0c"),u'(x"6c"),u'(x"01"),u'(x"6c"),u'(x"01"),u'(x"45"),u'(x"ff"),u'(x"60"),u'(x"10"),u'(x"01"),u'(x"01"),u'(x"a0"),u'(x"00"),
u'(x"02"),u'(x"65"),u'(x"00"),u'(x"eb"),u'(x"01"),u'(x"a0"),u'(x"00"),u'(x"02"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"eb"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"eb"),
u'(x"00"),u'(x"0a"),u'(x"eb"),u'(x"15"),u'(x"01"),u'(x"0a"),u'(x"20"),u'(x"01"),u'(x"02"),u'(x"a0"),u'(x"00"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"eb"),u'(x"01"),
u'(x"a0"),u'(x"00"),u'(x"87"),u'(x"a0"),u'(x"00"),u'(x"82"),u'(x"15"),u'(x"00"),u'(x"eb"),u'(x"09"),u'(x"ff"),u'(x"01"),u'(x"00"),u'(x"ad"),u'(x"eb"),u'(x"00"),
u'(x"02"),u'(x"a0"),u'(x"00"),u'(x"02"),u'(x"09"),u'(x"f3"),u'(x"01"),u'(x"a0"),u'(x"00"),u'(x"02"),u'(x"09"),u'(x"f3"),u'(x"01"),u'(x"a0"),u'(x"00"),u'(x"02"),
u'(x"09"),u'(x"f3"),u'(x"01"),u'(x"a0"),u'(x"00"),u'(x"02"),u'(x"09"),u'(x"f3"),u'(x"01"),u'(x"a0"),u'(x"00"),u'(x"02"),u'(x"09"),u'(x"f3"),u'(x"01"),u'(x"ad"),
u'(x"ea"),u'(x"00"),u'(x"02"),u'(x"90"),u'(x"ea"),u'(x"90"),u'(x"ea"),u'(x"01"),u'(x"ad"),u'(x"ea"),u'(x"00"),u'(x"02"),u'(x"90"),u'(x"ea"),u'(x"90"),u'(x"ea"),
u'(x"01"),u'(x"ad"),u'(x"ea"),u'(x"00"),u'(x"02"),u'(x"8b"),u'(x"ea"),u'(x"03"),u'(x"8b"),u'(x"ea"),u'(x"02"),u'(x"e5"),u'(x"00"),u'(x"90"),u'(x"ea"),u'(x"01"),
u'(x"e5"),u'(x"00"),u'(x"10"),u'(x"ea"),u'(x"9d"),u'(x"ea"),u'(x"10"),u'(x"ea"),u'(x"8a"),u'(x"ea"),u'(x"09"),u'(x"fb"),u'(x"01"),u'(x"15"),u'(x"00"),u'(x"ea"),
u'(x"00"),u'(x"a0"),u'(x"00"),u'(x"02"),u'(x"01"),u'(x"90"),u'(x"ea"),u'(x"10"),u'(x"45"),u'(x"ff"),u'(x"0c"),u'(x"1c"),u'(x"1b"),u'(x"20"),u'(x"00"),u'(x"86"),
u'(x"10"),u'(x"ea"),u'(x"01"),u'(x"09"),u'(x"15"),u'(x"00"),u'(x"ea"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ea"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ea"),u'(x"00"),
u'(x"15"),u'(x"00"),u'(x"ea"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ea"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ea"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ea"),u'(x"00"),
u'(x"15"),u'(x"00"),u'(x"ea"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ea"),u'(x"00"),u'(x"10"),u'(x"10"),u'(x"0a"),u'(x"15"),u'(x"90"),u'(x"15"),u'(x"98"),u'(x"10"),
u'(x"20"),u'(x"02"),u'(x"15"),u'(x"15"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"1d"),u'(x"e9"),u'(x"1d"),u'(x"e9"),u'(x"20"),u'(x"02"),u'(x"0a"),u'(x"01"),
u'(x"0a"),u'(x"e9"),u'(x"0a"),u'(x"20"),u'(x"00"),u'(x"87"),u'(x"0a"),u'(x"10"),u'(x"e9"),u'(x"65"),u'(x"00"),u'(x"92"),u'(x"45"),u'(x"ff"),u'(x"8b"),u'(x"e9"),
u'(x"03"),u'(x"2d"),u'(x"e9"),u'(x"00"),u'(x"86"),u'(x"8b"),u'(x"e9"),u'(x"02"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"02"),u'(x"8a"),u'(x"e9"),u'(x"15"),u'(x"00"),
u'(x"ff"),u'(x"00"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"1d"),u'(x"e9"),u'(x"1d"),u'(x"e9"),u'(x"20"),u'(x"02"),u'(x"0a"),u'(x"01"),u'(x"0a"),u'(x"20"),u'(x"00"),
u'(x"87"),u'(x"0a"),u'(x"10"),u'(x"e9"),u'(x"65"),u'(x"00"),u'(x"92"),u'(x"45"),u'(x"ff"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"a0"),u'(x"00"),u'(x"02"),
u'(x"8b"),u'(x"e9"),u'(x"02"),u'(x"8a"),u'(x"e9"),u'(x"01"),u'(x"8a"),u'(x"e9"),u'(x"01"),u'(x"a0"),u'(x"00"),u'(x"02"),u'(x"8a"),u'(x"e9"),u'(x"a0"),u'(x"00"),
u'(x"02"),u'(x"8a"),u'(x"e9"),u'(x"00"),u'(x"10"),u'(x"a0"),u'(x"00"),u'(x"02"),u'(x"8b"),u'(x"e9"),u'(x"02"),u'(x"95"),u'(x"00"),u'(x"e9"),u'(x"0a"),u'(x"01"),
u'(x"95"),u'(x"00"),u'(x"e9"),u'(x"0a"),u'(x"01"),u'(x"a0"),u'(x"00"),u'(x"02"),u'(x"95"),u'(x"00"),u'(x"e9"),u'(x"0a"),u'(x"01"),u'(x"a0"),u'(x"00"),u'(x"02"),
u'(x"95"),u'(x"00"),u'(x"e8"),u'(x"0a"),u'(x"01"),u'(x"a0"),u'(x"00"),u'(x"02"),u'(x"8b"),u'(x"e8"),u'(x"03"),u'(x"8a"),u'(x"e8"),u'(x"0a"),u'(x"01"),u'(x"95"),
u'(x"00"),u'(x"e8"),u'(x"0a"),u'(x"01"),u'(x"00"),u'(x"8b"),u'(x"e8"),u'(x"03"),u'(x"09"),u'(x"ff"),u'(x"8a"),u'(x"e8"),u'(x"8a"),u'(x"e8"),u'(x"0a"),u'(x"00"),
u'(x"a0"),u'(x"00"),u'(x"02"),u'(x"90"),u'(x"e8"),u'(x"0a"),u'(x"00"),u'(x"a0"),u'(x"00"),u'(x"02"),u'(x"90"),u'(x"e8"),u'(x"0a"),u'(x"00"),u'(x"8b"),u'(x"e8"),
u'(x"03"),u'(x"8b"),u'(x"e8"),u'(x"02"),u'(x"09"),u'(x"ff"),u'(x"8a"),u'(x"e8"),u'(x"0b"),u'(x"03"),u'(x"8a"),u'(x"e8"),u'(x"45"),u'(x"ff"),u'(x"9c"),u'(x"1e"),
u'(x"8b"),u'(x"03"),u'(x"01"),u'(x"a0"),u'(x"00"),u'(x"02"),u'(x"95"),u'(x"00"),u'(x"e8"),u'(x"01"),u'(x"a0"),u'(x"00"),u'(x"02"),u'(x"95"),u'(x"00"),u'(x"e8"),
u'(x"01"),u'(x"09"),u'(x"ff"),u'(x"0b"),u'(x"02"),u'(x"01"),u'(x"b5"),u'(x"00"),u'(x"02"),u'(x"45"),u'(x"ff"),u'(x"8b"),u'(x"e8"),u'(x"02"),u'(x"8b"),u'(x"e8"),
u'(x"02"),u'(x"01"),u'(x"8b"),u'(x"e8"),u'(x"02"),u'(x"8b"),u'(x"e8"),u'(x"02"),u'(x"9c"),u'(x"1d"),u'(x"01"),u'(x"9c"),u'(x"1e"),u'(x"8b"),u'(x"03"),u'(x"a0"),
u'(x"00"),u'(x"87"),u'(x"a0"),u'(x"00"),u'(x"82"),u'(x"e5"),u'(x"00"),u'(x"a0"),u'(x"00"),u'(x"02"),u'(x"8a"),u'(x"e7"),u'(x"01"),u'(x"a0"),u'(x"00"),u'(x"02"),
u'(x"8a"),u'(x"e7"),u'(x"8a"),u'(x"e7"),u'(x"01"),u'(x"01"),u'(x"a0"),u'(x"00"),u'(x"03"),u'(x"a0"),u'(x"00"),u'(x"87"),u'(x"a0"),u'(x"00"),u'(x"82"),u'(x"e5"),
u'(x"00"),u'(x"01"),u'(x"8b"),u'(x"e7"),u'(x"02"),u'(x"8b"),u'(x"e7"),u'(x"02"),u'(x"8b"),u'(x"e7"),u'(x"02"),u'(x"9c"),u'(x"1d"),u'(x"01"),u'(x"9c"),u'(x"1e"),
u'(x"45"),u'(x"ff"),u'(x"8b"),u'(x"03"),u'(x"01"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"0a"),u'(x"00"),u'(x"8b"),u'(x"ff"),u'(x"80"),u'(x"10"),u'(x"10"),u'(x"97"),
u'(x"ff"),u'(x"1d"),u'(x"e7"),u'(x"0a"),u'(x"20"),u'(x"00"),u'(x"87"),u'(x"0a"),u'(x"20"),u'(x"e7"),u'(x"03"),u'(x"0a"),u'(x"e7"),u'(x"10"),u'(x"e7"),u'(x"65"),
u'(x"00"),u'(x"90"),u'(x"2d"),u'(x"e6"),u'(x"00"),u'(x"87"),u'(x"8b"),u'(x"e6"),u'(x"02"),u'(x"8a"),u'(x"e6"),u'(x"15"),u'(x"00"),u'(x"09"),u'(x"00"),u'(x"15"),
u'(x"15"),u'(x"15"),u'(x"00"),u'(x"ff"),u'(x"00"),u'(x"8b"),u'(x"ff"),u'(x"80"),u'(x"90"),u'(x"ff"),u'(x"00"),u'(x"00"),u'(x"8b"),u'(x"d0"),u'(x"80"),u'(x"10"),
u'(x"10"),u'(x"1d"),u'(x"e6"),u'(x"1d"),u'(x"e6"),u'(x"0a"),u'(x"20"),u'(x"00"),u'(x"87"),u'(x"0a"),u'(x"20"),u'(x"03"),u'(x"10"),u'(x"e6"),u'(x"97"),u'(x"d0"),
u'(x"65"),u'(x"00"),u'(x"90"),u'(x"15"),u'(x"15"),u'(x"15"),u'(x"00"),u'(x"d0"),u'(x"00"),u'(x"65"),u'(x"6c"),u'(x"2c"),u'(x"77"),u'(x"72"),u'(x"64"),u'(x"20"),
u'(x"50"),u'(x"50"),u'(x"30"),u'(x"31"),u'(x"76"),u'(x"31"),u'(x"30"),u'(x"00"),u'(x"65"),u'(x"6c"),u'(x"2c"),u'(x"77"),u'(x"72"),u'(x"64"),u'(x"20"),u'(x"50"),
u'(x"50"),u'(x"30"),u'(x"31"),u'(x"76"),u'(x"31"),u'(x"35"),u'(x"00"),u'(x"15"),u'(x"15"),u'(x"15"),u'(x"15"),u'(x"16"),u'(x"16"),u'(x"16"),u'(x"17"),u'(x"17"),
u'(x"17"),u'(x"17"),u'(x"17"),u'(x"17"),u'(x"17"),u'(x"17"),u'(x"17"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"0c"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"08"),u'(x"0e"),u'(x"10"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"0b"),u'(x"0b"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"0b"),u'(x"0b"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"0b"),u'(x"0b"),u'(x"0b"),u'(x"00"),u'(x"00"),u'(x"0b"),u'(x"0b"),u'(x"0b"),u'(x"0b"),u'(x"0b"),u'(x"0b"),u'(x"0b"),u'(x"0b"),
u'(x"0c"),u'(x"0c"),u'(x"0c"),u'(x"00"),u'(x"0c"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"0c"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"0c"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"14"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"14"),u'(x"00"),u'(x"00"),u'(x"14"),
u'(x"14"),u'(x"14"),u'(x"14"),u'(x"14"),u'(x"15"),u'(x"15"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"15"),
u'(x"00"),u'(x"15"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"0c"),u'(x"0c"),u'(x"0c"),u'(x"0c"),u'(x"0d"),u'(x"12"),u'(x"12"),u'(x"12"),u'(x"0d"),
u'(x"12"),u'(x"0d"),u'(x"0d"),u'(x"0d"),u'(x"0e"),u'(x"12"),u'(x"12"),u'(x"0e"),u'(x"12"),u'(x"12"),u'(x"12"),u'(x"12"),u'(x"12"),u'(x"12"),u'(x"12"),u'(x"0e"),
u'(x"12"),u'(x"12"),u'(x"12"),u'(x"12"),u'(x"12"),u'(x"12"),u'(x"12"),u'(x"12"),u'(x"12"),u'(x"12"),u'(x"0e"),u'(x"12"),u'(x"12"),u'(x"0f"),u'(x"0f"),u'(x"0f"),
u'(x"12"),u'(x"12"),u'(x"12"),u'(x"0f"),u'(x"10"),u'(x"10"),u'(x"12"),u'(x"12"),u'(x"12"),u'(x"11"),u'(x"12"),u'(x"12"),u'(x"12"),u'(x"12"),u'(x"12"),u'(x"11"),
u'(x"12"),u'(x"12"),u'(x"12"),u'(x"12"),u'(x"12"),u'(x"12"),u'(x"12"),u'(x"80"),u'(x"80"),u'(x"81"),u'(x"81"),u'(x"82"),u'(x"83"),u'(x"83"),u'(x"84"),u'(x"85"),
u'(x"85"),u'(x"86"),u'(x"86"),u'(x"87"),u'(x"88"),u'(x"88"),u'(x"89"),u'(x"8a"),u'(x"8a"),u'(x"8b"),u'(x"8b"),u'(x"8c"),u'(x"8d"),u'(x"8d"),u'(x"8e"),u'(x"8f"),
u'(x"00"),u'(x"00"),u'(x"fd"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"09"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"71"),u'(x"00"),u'(x"00"),u'(x"73"),u'(x"77"),u'(x"00"),
u'(x"63"),u'(x"64"),u'(x"34"),u'(x"00"),u'(x"20"),u'(x"66"),u'(x"72"),u'(x"00"),u'(x"6e"),u'(x"68"),u'(x"79"),u'(x"00"),u'(x"00"),u'(x"6a"),u'(x"37"),u'(x"00"),
u'(x"2c"),u'(x"69"),u'(x"30"),u'(x"00"),u'(x"2e"),u'(x"6c"),u'(x"70"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"3d"),u'(x"00"),u'(x"00"),u'(x"5d"),u'(x"5c"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"f0"),u'(x"f3"),u'(x"00"),u'(x"00"),u'(x"ee"),u'(x"f4"),u'(x"f7"),u'(x"e9"),u'(x"ed"),u'(x"ec"),u'(x"f8"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"09"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"51"),u'(x"00"),u'(x"00"),u'(x"53"),u'(x"57"),u'(x"00"),
u'(x"43"),u'(x"44"),u'(x"24"),u'(x"00"),u'(x"20"),u'(x"46"),u'(x"52"),u'(x"00"),u'(x"4e"),u'(x"48"),u'(x"59"),u'(x"00"),u'(x"00"),u'(x"4a"),u'(x"26"),u'(x"00"),
u'(x"3c"),u'(x"49"),u'(x"29"),u'(x"00"),u'(x"3e"),u'(x"4c"),u'(x"50"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"2b"),u'(x"00"),u'(x"00"),u'(x"7d"),u'(x"7c"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"fc"),u'(x"e1"),u'(x"00"),u'(x"00"),u'(x"fb"),u'(x"00"),u'(x"e4"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"e6"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),
u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00"),u'(x"00") 
);

begin
   base_addr_match <= '1' when base_addr(17 downto 13) = bus_addr(17 downto 13) else '0';
   bus_addr_match <= base_addr_match;

   process(clk, base_addr_match)
   begin
      if clk = '1' and clk'event then
         bus_dati(7 downto 0) <= meme(conv_integer(bus_addr(12 downto 1)));
         bus_dati(15 downto 8) <= memo(conv_integer(bus_addr(12 downto 1)));
      end if;
   end process;

   process(clk, base_addr_match)
   begin
      if clk = '1' and clk'event then
         if base_addr_match = '1' and bus_control_dato = '1' and bus_addr(12 downto 9) = "0000" then       -- only 0..1000 writable
            if bus_control_datob = '0' or (bus_control_datob = '1' and bus_addr(0) = '0') then
               meme(conv_integer(bus_addr(12 downto 1))) <= bus_dato(7 downto 0);
            end if;
            if bus_control_datob = '0' or (bus_control_datob = '1' and bus_addr(0) = '1') then
               memo(conv_integer(bus_addr(12 downto 1))) <= bus_dato(15 downto 8);
            end if;
         end if;
      end if;
   end process;
end implementation;

